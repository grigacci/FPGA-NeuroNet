library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.CONFIG.ALL;
use ieee.float_pkg.all;
use work.bfloat_pkg.ALL;

package mulmat_soft_mem is
    type bias_array is array (0 to output_classes - 1) of f4; 
    type float_matrix is array (0 to number_of_neurons -1,0 to output_classes - 1)  of  f4;

    constant soft_bias : bias_array := 
    (to_f4(-0.875),to_f4(-0.875),to_f4(-0.875),to_f4(0.875),to_f4(0.875),to_f4(-0.875),to_f4(0.750),to_f4(-0.750),to_f4(0.875),to_f4(-0.8));
    
    constant soft_weights : float_matrix := 
    ((to_f4(0.125),to_f4(-0.875),to_f4(-0.750),to_f4(0.250),to_f4(0.500),to_f4(0.875),to_f4(-0.875),to_f4(0.875),to_f4(0.375),to_f4(0.500)),
(to_f4(-0.875),to_f4(0.625),to_f4(-0.875),to_f4(-0.875),to_f4(-0.875),to_f4(0.875),to_f4(0.875),to_f4(0.125),to_f4(-0.625),to_f4(-0.375)),
(to_f4(-0.125),to_f4(0.875),to_f4(0.875),to_f4(0.375),to_f4(0.375),to_f4(-0.875),to_f4(-0.500),to_f4(0.000),to_f4(0.750),to_f4(0.875)),
(to_f4(0.375),to_f4(-0.875),to_f4(-0.875),to_f4(-0.750),to_f4(0.625),to_f4(0.375),to_f4(0.500),to_f4(0.000),to_f4(0.875),to_f4(0.500)),
(to_f4(-0.875),to_f4(0.875),to_f4(0.875),to_f4(0.500),to_f4(-0.875),to_f4(0.000),to_f4(-0.875),to_f4(0.875),to_f4(-0.625),to_f4(-0.875)),
(to_f4(-0.875),to_f4(-0.875),to_f4(0.750),to_f4(0.000),to_f4(0.875),to_f4(0.125),to_f4(0.500),to_f4(-0.875),to_f4(0.625),to_f4(0.500)),
(to_f4(-0.625),to_f4(-0.250),to_f4(0.250),to_f4(0.875),to_f4(-0.500),to_f4(0.875),to_f4(-0.875),to_f4(-0.875),to_f4(-0.750),to_f4(0.250)),
(to_f4(-0.875),to_f4(-0.875),to_f4(-0.750),to_f4(-0.125),to_f4(-0.875),to_f4(0.875),to_f4(0.750),to_f4(-0.750),to_f4(0.625),to_f4(-0.250)),
(to_f4(-0.875),to_f4(0.375),to_f4(-0.875),to_f4(0.375),to_f4(0.875),to_f4(0.375),to_f4(-0.625),to_f4(0.000),to_f4(0.625),to_f4(0.750)),
(to_f4(0.000),to_f4(0.625),to_f4(-0.125),to_f4(0.875),to_f4(-0.875),to_f4(0.875),to_f4(-0.750),to_f4(-0.875),to_f4(-0.875),to_f4(-0.375)),
(to_f4(0.875),to_f4(0.500),to_f4(0.875),to_f4(-0.625),to_f4(-0.250),to_f4(-0.500),to_f4(0.875),to_f4(-0.875),to_f4(-0.375),to_f4(-0.750)),
(to_f4(0.375),to_f4(0.875),to_f4(0.500),to_f4(0.875),to_f4(-0.875),to_f4(-0.750),to_f4(-0.875),to_f4(-0.125),to_f4(-0.375),to_f4(0.750)),
(to_f4(0.750),to_f4(-0.875),to_f4(0.375),to_f4(0.875),to_f4(-0.875),to_f4(-0.375),to_f4(-0.875),to_f4(0.125),to_f4(0.875),to_f4(0.875)),
(to_f4(0.875),to_f4(0.000),to_f4(0.125),to_f4(-0.875),to_f4(-0.875),to_f4(0.750),to_f4(0.375),to_f4(-0.250),to_f4(0.875),to_f4(-0.875)),
(to_f4(0.125),to_f4(0.000),to_f4(-0.375),to_f4(0.500),to_f4(-0.875),to_f4(0.625),to_f4(0.875),to_f4(0.125),to_f4(0.125),to_f4(-0.875)),
(to_f4(0.875),to_f4(-0.875),to_f4(0.875),to_f4(0.875),to_f4(-0.875),to_f4(-0.875),to_f4(-0.750),to_f4(0.375),to_f4(0.500),to_f4(0.625)),
(to_f4(0.500),to_f4(0.500),to_f4(-0.125),to_f4(-0.875),to_f4(0.875),to_f4(0.250),to_f4(0.125),to_f4(0.875),to_f4(-0.625),to_f4(0.500)),
(to_f4(-0.875),to_f4(-0.250),to_f4(0.375),to_f4(0.000),to_f4(-0.250),to_f4(-0.875),to_f4(-0.125),to_f4(0.875),to_f4(-0.875),to_f4(0.000)),
(to_f4(0.500),to_f4(0.875),to_f4(0.625),to_f4(-0.250),to_f4(0.875),to_f4(-0.125),to_f4(0.125),to_f4(0.250),to_f4(-0.875),to_f4(-0.125)),
(to_f4(-0.125),to_f4(0.750),to_f4(0.875),to_f4(-0.125),to_f4(0.000),to_f4(0.000),to_f4(0.000),to_f4(0.125),to_f4(0.875),to_f4(-0.8)));
 
end mulmat_soft_mem;