library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.bfloat_pkg.ALL;

package input_data is
    type input_array is array(natural range<>, natural range<>) of bfloat16;

    constant input_image : input_array(27 downto 0,27 downto 0) := 
    ((to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(-0.00001),to_float(-0.00003),to_float(-0.00001),to_float(-0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(-0.00000),to_float(-0.00000),to_float(-0.00004),to_float(-0.00009),to_float(-0.00017),to_float(-0.00025),to_float(-0.00047),to_float(-0.00063),to_float(-0.00068),to_float(-0.00069),to_float(-0.00074),to_float(-0.00068),to_float(-0.00073),to_float(-0.00060),to_float(-0.00039),to_float(-0.00028),to_float(-0.00021),to_float(-0.00008),to_float(-0.00004),to_float(-0.00001),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(-0.00000),to_float(-0.00000),to_float(-0.00003),to_float(-0.00002),to_float(-0.00018),to_float(-0.00054),to_float(-0.00103),to_float(-0.00198),to_float(-0.00339),to_float(-0.00504),to_float(-0.00731),to_float(-0.00988),to_float(-0.01250),to_float(-0.01416),to_float(-0.01454),to_float(-0.01325),to_float(-0.01095),to_float(-0.00799),to_float(-0.00470),to_float(-0.00247),to_float(-0.00116),to_float(-0.00037),to_float(-0.00014),to_float(-0.00003),to_float(0.00000),to_float(0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(-0.00001),to_float(-0.00002),to_float(-0.00005),to_float(-0.00027),to_float(-0.00083),to_float(-0.00213),to_float(-0.00451),to_float(-0.00866),to_float(-0.01421),to_float(-0.02124),to_float(-0.02893),to_float(-0.03787),to_float(-0.04642),to_float(-0.05170),to_float(-0.05127),to_float(-0.04614),to_float(-0.03729),to_float(-0.02681),to_float(-0.01639),to_float(-0.00889),to_float(-0.00414),to_float(-0.00161),to_float(-0.00063),to_float(-0.00011),to_float(-0.00001),to_float(0.00000)),
    (to_float(0.00000),to_float(-0.00000),to_float(-0.00002),to_float(-0.00006),to_float(-0.00032),to_float(-0.00160),to_float(-0.00407),to_float(-0.00945),to_float(-0.01866),to_float(-0.03278),to_float(-0.05200),to_float(-0.07611),to_float(-0.10559),to_float(-0.13757),to_float(-0.16345),to_float(-0.17676),to_float(-0.17322),to_float(-0.15295),to_float(-0.12238),to_float(-0.08954),to_float(-0.05792),to_float(-0.03384),to_float(-0.01776),to_float(-0.00835),to_float(-0.00337),to_float(-0.00081),to_float(-0.00012),to_float(-0.00001)),
    (to_float(0.00000),to_float(0.00000),to_float(-0.00004),to_float(-0.00025),to_float(-0.00154),to_float(-0.00572),to_float(-0.01402),to_float(-0.02823),to_float(-0.05084),to_float(-0.08289),to_float(-0.12305),to_float(-0.17273),to_float(-0.23010),to_float(-0.28833),to_float(-0.33252),to_float(-0.35400),to_float(-0.34741),to_float(-0.31323),to_float(-0.25757),to_float(-0.19446),to_float(-0.13416),to_float(-0.08405),to_float(-0.04840),to_float(-0.02594),to_float(-0.01169),to_float(-0.00330),to_float(-0.00055),to_float(-0.00002)),
    (to_float(0.00000),to_float(-0.00000),to_float(-0.00011),to_float(-0.00086),to_float(-0.00437),to_float(-0.01285),to_float(-0.02905),to_float(-0.05569),to_float(-0.09430),to_float(-0.14563),to_float(-0.20752),to_float(-0.27710),to_float(-0.34863),to_float(-0.41504),to_float(-0.46289),to_float(-0.48486),to_float(-0.47534),to_float(-0.43774),to_float(-0.37549),to_float(-0.29370),to_float(-0.21106),to_float(-0.13794),to_float(-0.08197),to_float(-0.04471),to_float(-0.02104),to_float(-0.00725),to_float(-0.00146),to_float(-0.00012)),
    (to_float(-0.00000),to_float(-0.00008),to_float(-0.00042),to_float(-0.00233),to_float(-0.00903),to_float(-0.02316),to_float(0.27954),to_float(0.63477),to_float(0.47949),to_float(0.37939),to_float(-0.05371),to_float(-0.22705),to_float(-0.43579),to_float(-0.48828),to_float(-0.51855),to_float(-0.52881),to_float(-0.52100),to_float(-0.49487),to_float(-0.44360),to_float(-0.36621),to_float(-0.27246),to_float(-0.18298),to_float(-0.10992),to_float(-0.05939),to_float(-0.02748),to_float(-0.01009),to_float(-0.00200),to_float(-0.00012)),
    (to_float(-0.00002),to_float(-0.00020),to_float(-0.00129),to_float(-0.00515),to_float(-0.01464),to_float(-0.03314),to_float(0.80176),to_float(0.87646),to_float(0.80859),to_float(0.72607),to_float(0.63965),to_float(0.51758),to_float(0.30688),to_float(0.29150),to_float(0.29272),to_float(0.29565),to_float(0.29395),to_float(0.29639),to_float(0.31934),to_float(0.38037),to_float(0.36206),to_float(-0.00354),to_float(-0.12427),to_float(-0.06390),to_float(-0.02808),to_float(-0.01019),to_float(-0.00188),to_float(-0.00011)),
    (to_float(-0.00002),to_float(-0.00031),to_float(-0.00200),to_float(-0.00672),to_float(-0.01736),to_float(-0.03830),to_float(0.18542),to_float(0.31055),to_float(0.06763),to_float(0.14014),to_float(0.24976),to_float(0.45459),to_float(0.55957),to_float(0.47046),to_float(0.60547),to_float(0.60400),to_float(0.58496),to_float(0.54346),to_float(0.46069),to_float(0.60498),to_float(0.69141),to_float(0.34082),to_float(-0.12286),to_float(-0.06012),to_float(-0.02328),to_float(-0.00742),to_float(-0.00137),to_float(-0.00011)),
    (to_float(-0.00003),to_float(-0.00039),to_float(-0.00204),to_float(-0.00654),to_float(-0.01675),to_float(-0.03857),to_float(-0.08026),to_float(-0.14526),to_float(-0.23328),to_float(-0.32568),to_float(-0.39160),to_float(-0.33667),to_float(-0.10889),to_float(-0.26929),to_float(-0.04858),to_float(-0.06836),to_float(-0.10498),to_float(-0.17749),to_float(-0.33301),to_float(0.55371),to_float(0.71143),to_float(0.22534),to_float(-0.11127),to_float(-0.05273),to_float(-0.01797),to_float(-0.00449),to_float(-0.00087),to_float(-0.00007)),
    (to_float(-0.00002),to_float(-0.00030),to_float(-0.00164),to_float(-0.00500),to_float(-0.01424),to_float(-0.03732),to_float(-0.08258),to_float(-0.15564),to_float(-0.25024),to_float(-0.34058),to_float(-0.38574),to_float(-0.37061),to_float(-0.31909),to_float(-0.28638),to_float(-0.29736),to_float(-0.33374),to_float(-0.38013),to_float(-0.41992),to_float(-0.08789),to_float(0.64062),to_float(0.56250),to_float(-0.09570),to_float(-0.09900),to_float(-0.04913),to_float(-0.01559),to_float(-0.00236),to_float(-0.00049),to_float(-0.00003)),
    (to_float(-0.00001),to_float(-0.00017),to_float(-0.00095),to_float(-0.00343),to_float(-0.01199),to_float(-0.03754),to_float(-0.08899),to_float(-0.17017),to_float(-0.26953),to_float(-0.35254),to_float(-0.38232),to_float(-0.35571),to_float(-0.31128),to_float(-0.31006),to_float(-0.34888),to_float(-0.39722),to_float(-0.44165),to_float(-0.37329),to_float(0.49048),to_float(0.66602),to_float(0.09534),to_float(-0.14941),to_float(-0.09271),to_float(-0.04965),to_float(-0.01677),to_float(-0.00173),to_float(-0.00031),to_float(-0.00004)),
    (to_float(-0.00000),to_float(-0.00007),to_float(-0.00048),to_float(-0.00237),to_float(-0.01140),to_float(-0.04153),to_float(-0.09979),to_float(-0.18591),to_float(-0.28369),to_float(-0.35815),to_float(-0.37842),to_float(-0.35596),to_float(-0.33936),to_float(-0.37866),to_float(-0.43506),to_float(-0.48438),to_float(-0.50684),to_float(0.00928),to_float(0.56689),to_float(0.61230),to_float(-0.04382),to_float(-0.14539),to_float(-0.09363),to_float(-0.05328),to_float(-0.01993),to_float(-0.00228),to_float(-0.00032),to_float(-0.00004)),
    (to_float(-0.00001),to_float(-0.00003),to_float(-0.00021),to_float(-0.00182),to_float(-0.01198),to_float(-0.04825),to_float(-0.11145),to_float(-0.19727),to_float(-0.28809),to_float(-0.35303),to_float(-0.37134),to_float(-0.36450),to_float(-0.38208),to_float(-0.45093),to_float(-0.50879),to_float(-0.54492),to_float(-0.30518),to_float(0.47217),to_float(0.57422),to_float(-0.06860),to_float(-0.21912),to_float(-0.15210),to_float(-0.09973),to_float(-0.05710),to_float(-0.02235),to_float(-0.00320),to_float(-0.00036),to_float(-0.00001)),
    (to_float(-0.00000),to_float(-0.00002),to_float(-0.00018),to_float(-0.00197),to_float(-0.01391),to_float(-0.05627),to_float(-0.12103),to_float(-0.20007),to_float(-0.27905),to_float(-0.33496),to_float(-0.35693),to_float(-0.36816),to_float(-0.41040),to_float(-0.48120),to_float(-0.53027),to_float(-0.54346),to_float(0.00488),to_float(0.51758),to_float(0.33472),to_float(-0.28662),to_float(-0.22766),to_float(-0.16113),to_float(-0.10541),to_float(-0.05817),to_float(-0.02277),to_float(-0.00422),to_float(-0.00058),to_float(-0.00004)),
    (to_float(-0.00000),to_float(-0.00002),to_float(-0.00029),to_float(-0.00243),to_float(-0.01746),to_float(-0.06458),to_float(-0.12720),to_float(-0.19507),to_float(-0.25903),to_float(-0.30420),to_float(-0.32690),to_float(-0.34937),to_float(-0.39502),to_float(-0.45264),to_float(-0.49414),to_float(-0.46265),to_float(0.32788),to_float(0.53418),to_float(-0.14600),to_float(-0.30225),to_float(-0.23279),to_float(-0.16418),to_float(-0.10443),to_float(-0.05563),to_float(-0.02194),to_float(-0.00503),to_float(-0.00075),to_float(-0.00005)),
    (to_float(0.00000),to_float(-0.00003),to_float(-0.00044),to_float(-0.00372),to_float(-0.02325),to_float(-0.07239),to_float(-0.13062),to_float(-0.18823),to_float(-0.23621),to_float(-0.27026),to_float(-0.29175),to_float(-0.31543),to_float(-0.34985),to_float(-0.39819),to_float(-0.43994),to_float(0.04126),to_float(0.55371),to_float(0.30273),to_float(-0.36182),to_float(-0.30176),to_float(-0.23181),to_float(-0.15942),to_float(-0.09741),to_float(-0.05014),to_float(-0.02014),to_float(-0.00554),to_float(-0.00082),to_float(-0.00003)),
    (to_float(-0.00001),to_float(-0.00002),to_float(-0.00071),to_float(-0.00594),to_float(-0.02977),to_float(-0.07977),to_float(-0.13635),to_float(-0.18823),to_float(-0.22766),to_float(-0.25781),to_float(-0.28027),to_float(-0.29907),to_float(-0.32471),to_float(-0.37158),to_float(-0.12329),to_float(0.54199),to_float(0.50244),to_float(-0.18750),to_float(-0.36572),to_float(-0.29932),to_float(-0.22144),to_float(-0.14746),to_float(-0.08807),to_float(-0.04446),to_float(-0.01788),to_float(-0.00507),to_float(-0.00060),to_float(-0.00005)),
    (to_float(-0.00000),to_float(-0.00005),to_float(-0.00112),to_float(-0.00798),to_float(-0.03409),to_float(-0.08490),to_float(-0.14392),to_float(-0.19910),to_float(-0.24353),to_float(-0.27832),to_float(-0.30420),to_float(-0.32275),to_float(-0.35132),to_float(-0.32202),to_float(0.42407),to_float(0.53223),to_float(0.19556),to_float(-0.41968),to_float(-0.36035),to_float(-0.28076),to_float(-0.19849),to_float(-0.12769),to_float(-0.07330),to_float(-0.03577),to_float(-0.01422),to_float(-0.00417),to_float(-0.00057),to_float(-0.00003)),
    (to_float(0.00000),to_float(-0.00006),to_float(-0.00130),to_float(-0.00881),to_float(-0.03326),to_float(-0.08081),to_float(-0.14490),to_float(-0.21008),to_float(-0.26904),to_float(-0.31714),to_float(-0.35303),to_float(-0.38232),to_float(-0.40527),to_float(0.33472),to_float(0.50391),to_float(0.36499),to_float(-0.32495),to_float(-0.40552),to_float(-0.32764),to_float(-0.23926),to_float(-0.15991),to_float(-0.09741),to_float(-0.05322),to_float(-0.02554),to_float(-0.01060),to_float(-0.00293),to_float(-0.00044),to_float(-0.00001)),
    (to_float(-0.00000),to_float(-0.00005),to_float(-0.00111),to_float(-0.00718),to_float(-0.02591),to_float(-0.06604),to_float(-0.12817),to_float(-0.20142),to_float(-0.27515),to_float(-0.34082),to_float(-0.39453),to_float(-0.43921),to_float(-0.33057),to_float(0.48291),to_float(0.47705),to_float(-0.18701),to_float(-0.42969),to_float(-0.34937),to_float(-0.26001),to_float(-0.17810),to_float(-0.11157),to_float(-0.06366),to_float(-0.03323),to_float(-0.01605),to_float(-0.00665),to_float(-0.00173),to_float(-0.00023),to_float(-0.00000)),
    (to_float(-0.00000),to_float(-0.00000),to_float(-0.00073),to_float(-0.00425),to_float(-0.01541),to_float(-0.04236),to_float(-0.09137),to_float(-0.15869),to_float(-0.23816),to_float(-0.31641),to_float(-0.38721),to_float(-0.32080),to_float(0.39648),to_float(0.50293),to_float(-0.02197),to_float(-0.41479),to_float(-0.34253),to_float(-0.25781),to_float(-0.17712),to_float(-0.11224),to_float(-0.06604),to_float(-0.03580),to_float(-0.01839),to_float(-0.00869),to_float(-0.00326),to_float(-0.00074),to_float(-0.00007),to_float(-0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(-0.00025),to_float(-0.00164),to_float(-0.00677),to_float(-0.01959),to_float(-0.04700),to_float(-0.09351),to_float(-0.15723),to_float(-0.23010),to_float(-0.30176),to_float(0.15991),to_float(0.60254),to_float(0.60449),to_float(-0.15063),to_float(-0.29517),to_float(-0.22498),to_float(-0.15698),to_float(-0.09961),to_float(-0.05954),to_float(-0.03329),to_float(-0.01726),to_float(-0.00861),to_float(-0.00383),to_float(-0.00121),to_float(-0.00023),to_float(-0.00004),to_float(0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(-0.00006),to_float(-0.00048),to_float(-0.00212),to_float(-0.00625),to_float(-0.01642),to_float(-0.03571),to_float(-0.06573),to_float(-0.10577),to_float(0.08948),to_float(0.76172),to_float(0.79053),to_float(0.79297),to_float(0.02563),to_float(-0.14355),to_float(-0.10718),to_float(-0.07465),to_float(-0.04733),to_float(-0.02818),to_float(-0.01546),to_float(-0.00779),to_float(-0.00372),to_float(-0.00156),to_float(-0.00040),to_float(-0.00009),to_float(-0.00001),to_float(0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(-0.00001),to_float(-0.00007),to_float(-0.00050),to_float(-0.00185),to_float(-0.00549),to_float(-0.01243),to_float(-0.02400),to_float(-0.03839),to_float(0.41846),to_float(0.92676),to_float(0.92139),to_float(0.78613),to_float(0.09448),to_float(-0.05127),to_float(-0.04102),to_float(-0.03044),to_float(-0.02040),to_float(-0.01235),to_float(-0.00661),to_float(-0.00322),to_float(-0.00145),to_float(-0.00055),to_float(-0.00012),to_float(-0.00001),to_float(-0.00001),to_float(0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(-0.00000),to_float(-0.00014),to_float(-0.00064),to_float(-0.00210),to_float(-0.00468),to_float(-0.00905),to_float(-0.01372),to_float(0.45361),to_float(0.96875),to_float(0.78320),to_float(0.04587),to_float(-0.02176),to_float(-0.01738),to_float(-0.01381),to_float(-0.01012),to_float(-0.00665),to_float(-0.00394),to_float(-0.00211),to_float(-0.00093),to_float(-0.00029),to_float(-0.00006),to_float(-0.00000),to_float(-0.00000),to_float(0.00000),to_float(0.00000)),
    (to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(-0.00001),to_float(-0.00006),to_float(-0.00016),to_float(-0.00035),to_float(-0.00050),to_float(-0.00077),to_float(-0.00131),to_float(-0.00168),to_float(-0.00205),to_float(-0.00231),to_float(-0.00269),to_float(-0.00231),to_float(-0.00189),to_float(-0.00134),to_float(-0.00078),to_float(-0.00035),to_float(-0.00018),to_float(-0.00008),to_float(-0.00006),to_float(-0.00001),to_float(0.00000),to_float(0.00000),to_float(0.00000),to_float(0.00000)));

end package;    