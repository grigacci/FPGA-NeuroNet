library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.CONFIG.ALL;
use ieee.float_pkg.all;

package mulmat_mem is
    type float_matrix is array (0 to number_of_neurons - 1,0 to input_size -1)  of  float(weight_size/2 downto -weight_size/2);
    constant weights : float_matrix := 
    ((to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000)),
    (to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125)),
    (to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(0.250),to_float(0.125),to_float(-0.875),to_float(-0.375),to_float(0.250),to_float(0.500),to_float(0.875),to_float(-0.250),to_float(0.125),to_float(0.250)),
    (to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(-0.625),to_float(0.875),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(0.375),to_float(-0.875),to_float(0.250),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(0.250),to_float(0.875)),
    (to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.250),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.250),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(0.750),to_float(0.125),to_float(0.875),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.875)),
    (to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(0.625),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.250)),
    (to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000)),
    (to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125)),
    (to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.375),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.125)),
    (to_float(-0.125),to_float(-0.750),to_float(-0.500),to_float(0.625),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(-0.625),to_float(0.125),to_float(0.250),to_float(0.750),to_float(-0.125),to_float(0.125),to_float(0.125)),
    (to_float(-0.625),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.000),to_float(0.875),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(-0.625),to_float(0.375),to_float(-0.875),to_float(-0.625),to_float(0.250),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(0.000)),
    (to_float(-0.500),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.125),to_float(0.875),to_float(0.000),to_float(-0.375),to_float(-0.750),to_float(-0.375),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(0.000)),
    (to_float(-0.375),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.750),to_float(0.125),to_float(0.875),to_float(-0.375),to_float(-0.375),to_float(-0.375),to_float(0.000),to_float(-0.625),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(-0.375),to_float(0.875),to_float(0.000),to_float(0.250),to_float(0.500)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.500),to_float(0.250),to_float(0.875),to_float(0.000),to_float(-0.125),to_float(-0.500),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(0.250),to_float(0.875),to_float(0.125),to_float(0.375),to_float(0.250)),
    (to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.125),to_float(0.875),to_float(0.375),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(-0.250),to_float(0.875),to_float(-0.125),to_float(0.250),to_float(0.250)),
    (to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(0.750),to_float(-0.375),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(0.250),to_float(0.875)),
    (to_float(0.250),to_float(0.875),to_float(0.375),to_float(0.875),to_float(0.000),to_float(0.000),to_float(0.875),to_float(-0.375),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(0.875)),
    (to_float(0.500),to_float(0.500),to_float(-0.125),to_float(0.875),to_float(0.250),to_float(0.250),to_float(0.875),to_float(-0.750),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(-0.875)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.500),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.750),to_float(0.875),to_float(0.875),to_float(0.250),to_float(-0.875)),
    (to_float(-0.875),to_float(0.375),to_float(0.125),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.750),to_float(0.500),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.500),to_float(0.000),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.875)),
    (to_float(-0.750),to_float(-0.625),to_float(0.625),to_float(0.500),to_float(-0.250),to_float(0.125),to_float(0.750),to_float(0.375),to_float(-0.125),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(-0.375),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(0.500),to_float(-0.125),to_float(-0.375),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(-0.125),to_float(0.875),to_float(-0.375),to_float(-0.250),to_float(-0.250)),
    (to_float(-0.625),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.750),to_float(-0.250),to_float(0.875),to_float(0.625),to_float(-0.500),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(0.625),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.500)),
    (to_float(-0.750),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.750),to_float(-0.250),to_float(0.875),to_float(0.500),to_float(-0.375),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.625)),
    (to_float(-0.750),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.250),to_float(-0.250),to_float(0.875),to_float(0.625),to_float(-0.375),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.000),to_float(0.875),to_float(-0.750),to_float(0.000),to_float(0.625)),
    (to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.125),to_float(0.875),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.500)),
    (to_float(-0.750),to_float(-0.250),to_float(-0.375),to_float(0.875),to_float(0.375),to_float(0.125),to_float(0.875),to_float(0.750),to_float(-0.125),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.250),to_float(0.500),to_float(0.875),to_float(-0.625),to_float(-0.625),to_float(0.250)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125)),
    (to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.000)),
    (to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.250),to_float(-0.125),to_float(0.750),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(0.875),to_float(-0.625),to_float(-0.125),to_float(0.000)),
    (to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.500),to_float(0.375),to_float(0.000),to_float(-0.625),to_float(-0.375),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.375),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(0.125),to_float(0.875),to_float(0.000),to_float(-0.625),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.875)),
    (to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.125),to_float(0.875),to_float(0.250),to_float(-0.500),to_float(-0.250),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.125),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(0.125)),
    (to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.375),to_float(0.875),to_float(0.000),to_float(-0.750),to_float(-0.625),to_float(0.375),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(-0.750),to_float(0.875),to_float(-0.375),to_float(0.000),to_float(0.500)),
    (to_float(-0.250),to_float(0.000),to_float(0.625),to_float(0.875),to_float(0.750),to_float(-0.375),to_float(0.875),to_float(-0.625),to_float(-0.875),to_float(-0.875),to_float(-0.625),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.875)),
    (to_float(0.500),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(0.125),to_float(0.250),to_float(-0.375),to_float(0.500),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.125),to_float(0.500),to_float(0.875)),
    (to_float(0.375),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(0.125),to_float(-0.125)),
    (to_float(-0.250),to_float(0.500),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(-0.750),to_float(0.875),to_float(0.375),to_float(-0.125),to_float(-0.750),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(-0.875)),
    (to_float(0.875),to_float(0.625),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.000),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.125),to_float(0.875),to_float(-0.250),to_float(-0.125),to_float(0.875),to_float(-0.375),to_float(-0.750),to_float(0.750)),
    (to_float(0.625),to_float(-0.500),to_float(0.750),to_float(0.750),to_float(-0.625),to_float(-0.125),to_float(-0.500),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(-0.625),to_float(-0.250),to_float(0.875),to_float(-0.375),to_float(0.000),to_float(-0.875),to_float(0.875)),
    (to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(-0.250),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(-0.875)),
    (to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(-0.500),to_float(0.875),to_float(-0.875),to_float(-0.875)),
    (to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.125),to_float(-0.625)),
    (to_float(-0.625),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.375),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(-0.750),to_float(-0.625),to_float(-0.625),to_float(0.625),to_float(0.875)),
    (to_float(-0.875),to_float(0.375),to_float(-0.125),to_float(0.875),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(0.875),to_float(0.750),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(0.875)),
    (to_float(0.750),to_float(0.875),to_float(0.000),to_float(0.875),to_float(-0.500),to_float(0.375),to_float(0.875),to_float(0.250),to_float(0.875),to_float(-0.125),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.875),to_float(-0.750),to_float(-0.125),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(-0.375),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.875)),
    (to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(0.500),to_float(-0.500),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(-0.625),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(0.875)),
    (to_float(-0.875),to_float(0.750),to_float(0.375),to_float(0.625),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.250),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.750),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(0.125)),
    (to_float(-0.875),to_float(-0.750),to_float(-0.125),to_float(0.875),to_float(0.250),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(-0.500),to_float(-0.250),to_float(0.875),to_float(-0.250),to_float(-0.625),to_float(-0.500)),
    (to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.750),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.375),to_float(-0.250),to_float(0.875),to_float(0.625),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.500),to_float(0.625),to_float(-0.250),to_float(-0.875),to_float(0.875)),
    (to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.250),to_float(-0.125),to_float(-0.625),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(-0.500),to_float(-0.375),to_float(-0.875),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(0.875),to_float(0.625),to_float(-0.375),to_float(-0.250)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125)),
    (to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(-0.250),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.125)),
    (to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(-0.375),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.250)),
    (to_float(0.000),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(0.125),to_float(0.750)),
    (to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(0.250),to_float(-0.875)),
    (to_float(0.000),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(0.375),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.625),to_float(0.125),to_float(0.625),to_float(-0.875)),
    (to_float(0.375),to_float(0.625),to_float(0.750),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(-0.875)),
    (to_float(0.625),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(0.375),to_float(-0.375),to_float(0.875),to_float(0.750),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(-0.375),to_float(0.875),to_float(0.500),to_float(0.500),to_float(-0.375),to_float(0.500),to_float(0.875)),
    (to_float(0.125),to_float(0.125),to_float(0.375),to_float(0.750),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(-0.500),to_float(-0.125),to_float(-0.875),to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(-0.375),to_float(0.875),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(0.875)),
    (to_float(0.875),to_float(-0.500),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(-0.125),to_float(0.750),to_float(0.750),to_float(0.250)),
    (to_float(0.875),to_float(-0.625),to_float(0.875),to_float(0.625),to_float(0.750),to_float(0.375),to_float(-0.875),to_float(0.375),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(-0.375),to_float(0.625),to_float(0.875),to_float(-0.625)),
    (to_float(0.500),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(-0.625),to_float(0.500),to_float(0.125),to_float(0.500),to_float(0.125),to_float(-0.625),to_float(-0.250),to_float(0.625)),
    (to_float(0.625),to_float(-0.125),to_float(0.625),to_float(0.125),to_float(0.625),to_float(0.375),to_float(0.625),to_float(-0.500),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(-0.750),to_float(0.375),to_float(-0.500),to_float(0.375),to_float(0.500),to_float(-0.375),to_float(-0.875),to_float(0.625)),
    (to_float(0.375),to_float(-0.625),to_float(0.875),to_float(0.625),to_float(0.250),to_float(0.625),to_float(-0.375),to_float(0.000),to_float(0.750),to_float(-0.750),to_float(-0.875),to_float(-0.625),to_float(-0.125),to_float(0.625),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.625),to_float(-0.375)),
    (to_float(-0.750),to_float(0.000),to_float(0.375),to_float(0.500),to_float(0.875),to_float(0.375),to_float(0.375),to_float(0.250),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.000),to_float(-0.625),to_float(0.000),to_float(-0.875),to_float(0.375),to_float(-0.625),to_float(0.125)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.625),to_float(-0.625),to_float(0.875),to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(-0.250),to_float(0.125),to_float(0.375),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(0.375)),
    (to_float(-0.875),to_float(-0.625),to_float(0.125),to_float(0.000),to_float(0.875),to_float(-0.750),to_float(0.500),to_float(-0.875),to_float(0.125),to_float(0.500),to_float(-0.875),to_float(0.250),to_float(0.250),to_float(0.500),to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.625)),
    (to_float(-0.500),to_float(0.375),to_float(0.000),to_float(0.500),to_float(0.250),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(-0.875)),
    (to_float(0.250),to_float(-0.875),to_float(-0.125),to_float(0.750),to_float(0.875),to_float(0.875),to_float(0.000),to_float(-0.125),to_float(0.750),to_float(-0.375),to_float(-0.750),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(0.625),to_float(-0.750),to_float(-0.875),to_float(-0.875)),
    (to_float(0.000),to_float(-0.250),to_float(0.750),to_float(0.625),to_float(-0.250),to_float(0.125),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.500),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.125),to_float(0.500)),
    (to_float(-0.250),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.500),to_float(-0.375),to_float(-0.625),to_float(0.375),to_float(0.375),to_float(0.000),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.125),to_float(0.375),to_float(0.875),to_float(0.625),to_float(0.500)),
    (to_float(0.875),to_float(-0.625),to_float(0.875),to_float(-0.250),to_float(0.375),to_float(0.875),to_float(0.625),to_float(-0.125),to_float(-0.875),to_float(-0.500),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.250),to_float(0.875)),
    (to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875)),
    (to_float(-0.125),to_float(-0.500),to_float(-0.500),to_float(0.875),to_float(0.625),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(-0.500),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.875)),
    (to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.500),to_float(0.875),to_float(0.250),to_float(0.000),to_float(0.875),to_float(-0.125)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125)),
    (to_float(0.000),to_float(-0.625),to_float(-0.375),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.750),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(0.625),to_float(-0.125),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(-0.875),to_float(0.750),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(-0.125),to_float(0.125),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.125)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(0.750),to_float(0.750),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.250)),
    (to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(0.750),to_float(0.875),to_float(-0.375),to_float(-0.750),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.375),to_float(0.500),to_float(0.875),to_float(0.250),to_float(-0.250),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.375),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.125)),
    (to_float(-0.875),to_float(0.750),to_float(0.750),to_float(-0.750),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.125)),
    (to_float(0.875),to_float(-0.625),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.625),to_float(-0.500),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(-0.875)),
    (to_float(-0.500),to_float(-0.375),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(0.375),to_float(-0.500),to_float(-0.625),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(0.250)),
    (to_float(0.125),to_float(0.625),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(0.750),to_float(-0.625),to_float(-0.500),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(-0.500),to_float(-0.125),to_float(0.250)),
    (to_float(0.000),to_float(0.625),to_float(0.750),to_float(0.125),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.125),to_float(-0.250),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.750),to_float(-0.875),to_float(0.750),to_float(0.500),to_float(0.375),to_float(-0.875),to_float(0.125)),
    (to_float(0.500),to_float(0.125),to_float(0.375),to_float(0.625),to_float(-0.625),to_float(0.875),to_float(-0.250),to_float(-0.375),to_float(0.500),to_float(-0.500),to_float(-0.250),to_float(-0.250),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(0.625),to_float(-0.750),to_float(0.500)),
    (to_float(0.500),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(-0.250),to_float(0.750),to_float(-0.375),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.125),to_float(0.750),to_float(0.625),to_float(-0.625),to_float(0.250),to_float(0.500),to_float(0.125),to_float(-0.875),to_float(-0.250)),
    (to_float(-0.375),to_float(-0.500),to_float(0.625),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(-0.750),to_float(0.250),to_float(-0.250),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(-0.125)),
    (to_float(0.500),to_float(-0.375),to_float(-0.125),to_float(0.625),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(-0.750),to_float(-0.875),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(0.000),to_float(0.375),to_float(-0.625),to_float(-0.500),to_float(-0.625),to_float(0.125)),
    (to_float(-0.125),to_float(0.125),to_float(-0.250),to_float(0.625),to_float(-0.250),to_float(0.625),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.625),to_float(-0.875),to_float(-0.125),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(0.625),to_float(0.375),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(0.125),to_float(0.375),to_float(-0.750),to_float(-0.125),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(0.000)),
    (to_float(-0.125),to_float(0.500),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(-0.250),to_float(0.125),to_float(-0.500),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(0.125),to_float(0.875),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(0.375)),
    (to_float(-0.625),to_float(-0.375),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.500),to_float(-0.500),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(0.375),to_float(0.375),to_float(-0.625),to_float(-0.125),to_float(0.750),to_float(-0.375)),
    (to_float(-0.125),to_float(0.125),to_float(0.625),to_float(0.750),to_float(-0.125),to_float(0.250),to_float(0.750),to_float(0.375),to_float(-0.250),to_float(0.125),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.250),to_float(0.875),to_float(0.000),to_float(-0.125),to_float(-0.250)),
    (to_float(0.500),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.500),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(0.375),to_float(0.000),to_float(-0.375),to_float(0.750),to_float(0.875),to_float(0.000),to_float(-0.500),to_float(0.500)),
    (to_float(-0.625),to_float(0.000),to_float(0.500),to_float(0.375),to_float(0.750),to_float(-0.375),to_float(0.250),to_float(0.500),to_float(-0.875),to_float(-0.125),to_float(0.625),to_float(0.125),to_float(-0.125),to_float(-0.500),to_float(0.000),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(0.875),to_float(-0.375)),
    (to_float(-0.625),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.125),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(-0.625),to_float(-0.500),to_float(-0.250),to_float(-0.625),to_float(-0.375),to_float(0.125)),
    (to_float(0.750),to_float(-0.750),to_float(-0.375),to_float(0.500),to_float(0.250),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(-0.625),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(-0.125)),
    (to_float(0.875),to_float(0.250),to_float(-0.875),to_float(0.250),to_float(-0.625),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.125),to_float(0.375),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(-0.875)),
    (to_float(0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.625),to_float(-0.625),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875)),
    (to_float(0.375),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.125),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.375),to_float(-0.500),to_float(0.500),to_float(-0.875)),
    (to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.250),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.625)),
    (to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.875)),
    (to_float(-0.250),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(0.250),to_float(0.500),to_float(-0.875),to_float(0.500),to_float(-0.375),to_float(-0.625),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(0.500),to_float(-0.750),to_float(0.125),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.375),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(0.750),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.250),to_float(0.750),to_float(-0.375),to_float(-0.875)),
    (to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.125),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.250),to_float(0.875),to_float(-0.625),to_float(0.875),to_float(-0.750)),
    (to_float(-0.875),to_float(-0.500),to_float(0.625),to_float(0.125),to_float(0.500),to_float(0.000),to_float(-0.625),to_float(0.875),to_float(0.000),to_float(-0.500),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(-0.750),to_float(0.500),to_float(-0.375),to_float(0.750),to_float(0.750),to_float(-0.125),to_float(0.125)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(-0.125),to_float(0.500),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(0.375),to_float(0.750),to_float(-0.625),to_float(0.375),to_float(-0.125)),
    (to_float(-0.250),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(-0.750),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(0.000),to_float(-0.375),to_float(-0.500),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.375),to_float(-0.750),to_float(0.250)),
    (to_float(-0.125),to_float(0.500),to_float(-0.500),to_float(0.375),to_float(0.250),to_float(-0.250),to_float(0.625),to_float(-0.625),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.500),to_float(0.375),to_float(0.750),to_float(0.000),to_float(-0.875),to_float(0.250)),
    (to_float(0.125),to_float(-0.250),to_float(0.375),to_float(0.125),to_float(0.250),to_float(0.500),to_float(0.250),to_float(-0.125),to_float(0.000),to_float(-0.625),to_float(0.500),to_float(0.125),to_float(0.000),to_float(-0.750),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.125),to_float(-0.875),to_float(0.375)),
    (to_float(0.000),to_float(-0.750),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(0.125),to_float(0.250),to_float(0.125),to_float(0.500),to_float(0.625),to_float(-0.125),to_float(-0.125),to_float(0.625),to_float(-0.375),to_float(-0.125),to_float(0.125),to_float(-0.750),to_float(-0.375),to_float(-0.250),to_float(0.250)),
    (to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.750),to_float(0.750),to_float(0.250),to_float(-0.250),to_float(0.250),to_float(-0.250),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(-0.625),to_float(-0.750),to_float(-0.250)),
    (to_float(-0.875),to_float(0.125),to_float(-0.500),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.500),to_float(-0.250),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(0.000),to_float(-0.625),to_float(0.000),to_float(-0.875),to_float(0.875)),
    (to_float(0.250),to_float(-0.125),to_float(0.625),to_float(0.125),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.500),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.375),to_float(-0.375),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(-0.625),to_float(-0.125)),
    (to_float(-0.875),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.375),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.125),to_float(-0.750),to_float(-0.375),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.500)),
    (to_float(0.125),to_float(-0.500),to_float(0.000),to_float(-0.375),to_float(0.000),to_float(0.500),to_float(0.250),to_float(-0.375),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(0.375),to_float(-0.250),to_float(0.375),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.000)),
    (to_float(0.250),to_float(-0.625),to_float(-0.375),to_float(0.625),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(-0.500),to_float(-0.125),to_float(0.500),to_float(-0.250),to_float(-0.375),to_float(0.250),to_float(-0.125),to_float(0.625),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(-0.750),to_float(-0.125)),
    (to_float(-0.625),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(0.375),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(-0.250),to_float(0.375),to_float(-0.250),to_float(-0.750),to_float(0.500),to_float(-0.250),to_float(0.250),to_float(-0.625),to_float(0.125)),
    (to_float(0.625),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(-0.250),to_float(0.625),to_float(-0.500),to_float(-0.625),to_float(0.500),to_float(-0.875),to_float(0.125),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(-0.375),to_float(-0.250),to_float(-0.250),to_float(-0.500),to_float(0.250),to_float(0.250)),
    (to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.375),to_float(0.875),to_float(-0.750),to_float(0.500),to_float(-0.625),to_float(-0.500),to_float(-0.500),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(0.625),to_float(0.500),to_float(0.000),to_float(-0.250)),
    (to_float(0.500),to_float(0.125),to_float(-0.500),to_float(0.375),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.625),to_float(0.500),to_float(0.000),to_float(0.625),to_float(0.250),to_float(0.500),to_float(0.625),to_float(-0.375),to_float(-0.625),to_float(0.375),to_float(-0.250),to_float(-0.750),to_float(-0.375)),
    (to_float(0.375),to_float(-0.500),to_float(-0.500),to_float(0.750),to_float(-0.625),to_float(-0.125),to_float(0.375),to_float(-0.875),to_float(0.750),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.375),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(-0.625),to_float(-0.500),to_float(0.125)),
    (to_float(-0.875),to_float(-0.750),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(0.125),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(-0.125),to_float(-0.375),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(-0.375),to_float(-0.875)),
    (to_float(0.000),to_float(-0.125),to_float(-0.375),to_float(-0.625),to_float(-0.500),to_float(0.000),to_float(-0.125),to_float(-0.625),to_float(-0.875),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.125),to_float(-0.750),to_float(0.375),to_float(-0.375),to_float(-0.375),to_float(-0.250)),
    (to_float(0.875),to_float(0.625),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(-0.625),to_float(0.000),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(-0.625)),
    (to_float(-0.125),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.750),to_float(0.125),to_float(0.625),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.000),to_float(-0.750),to_float(0.250),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(-0.625),to_float(0.750)),
    (to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.625),to_float(-0.375),to_float(-0.375),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.125)),
    (to_float(0.000),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(0.250),to_float(0.000),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(0.500),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.375)),
    (to_float(0.875),to_float(0.250),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.625),to_float(0.750),to_float(0.125),to_float(-0.250)),
    (to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(-0.250),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.375),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.625),to_float(-0.750),to_float(-0.500),to_float(-0.375)),
    (to_float(-0.500),to_float(0.375),to_float(0.875),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(0.875),to_float(-0.875)),
    (to_float(0.500),to_float(0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.625),to_float(-0.375),to_float(-0.875),to_float(0.750),to_float(0.750),to_float(0.750),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.250)),
    (to_float(0.000),to_float(0.125),to_float(-0.250),to_float(-0.750),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(0.875),to_float(0.000),to_float(-0.750),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.125),to_float(-0.625)),
    (to_float(0.250),to_float(-0.250),to_float(0.000),to_float(-0.375),to_float(-0.625),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(-0.625),to_float(-0.500),to_float(-0.625),to_float(-0.375),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.375)),
    (to_float(0.125),to_float(0.250),to_float(-0.625),to_float(0.000),to_float(0.500),to_float(0.250),to_float(0.250),to_float(0.250),to_float(-0.625),to_float(-0.250),to_float(0.500),to_float(0.000),to_float(-0.125),to_float(-0.625),to_float(-0.625),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(-0.250),to_float(0.000)),
    (to_float(-0.125),to_float(0.750),to_float(-0.625),to_float(-0.375),to_float(0.250),to_float(0.500),to_float(-0.375),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(-0.500),to_float(0.750),to_float(-0.875)),
    (to_float(-0.375),to_float(-0.125),to_float(0.500),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.625),to_float(-0.375),to_float(-0.500),to_float(0.125),to_float(0.375),to_float(0.125),to_float(0.625),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(0.250)),
    (to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.750),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(0.625),to_float(0.625),to_float(-0.250),to_float(-0.500),to_float(-0.125),to_float(0.375)),
    (to_float(0.000),to_float(0.500),to_float(-0.250),to_float(0.250),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.125),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(0.250),to_float(-0.500),to_float(-0.250),to_float(-0.375),to_float(0.125)),
    (to_float(-0.625),to_float(0.125),to_float(0.375),to_float(0.375),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(-0.250)),
    (to_float(0.375),to_float(-0.250),to_float(-0.500),to_float(0.625),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(0.750),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(-0.875),to_float(-0.500),to_float(-0.250),to_float(0.250)),
    (to_float(-0.750),to_float(-0.250),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.500),to_float(-0.250),to_float(-0.750),to_float(-0.250),to_float(0.000),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(0.625),to_float(0.000)),
    (to_float(-0.875),to_float(0.375),to_float(0.000),to_float(0.625),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(-0.375),to_float(-0.250),to_float(0.000),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(-0.250),to_float(0.625)),
    (to_float(0.125),to_float(0.500),to_float(-0.500),to_float(0.500),to_float(0.500),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(0.250),to_float(-0.750),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.500),to_float(0.125),to_float(0.125)),
    (to_float(-0.375),to_float(-0.125),to_float(-0.500),to_float(0.750),to_float(0.875),to_float(-0.125),to_float(-0.250),to_float(0.375),to_float(0.125),to_float(0.500),to_float(-0.125),to_float(-0.625),to_float(0.000),to_float(-0.125),to_float(-0.375),to_float(-0.375),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.500)),
    (to_float(0.375),to_float(0.000),to_float(-0.375),to_float(0.625),to_float(0.250),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.000),to_float(-0.625),to_float(-0.500),to_float(0.000),to_float(0.000),to_float(0.375),to_float(0.125),to_float(-0.125),to_float(-0.500),to_float(0.500)),
    (to_float(0.000),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.250),to_float(-0.750),to_float(0.125),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.375),to_float(-0.750),to_float(0.000),to_float(0.500),to_float(0.000),to_float(-0.375),to_float(0.250)),
    (to_float(-0.875),to_float(0.500),to_float(0.000),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(-0.750),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(0.125),to_float(0.125)),
    (to_float(0.375),to_float(-0.625),to_float(0.500),to_float(-0.875),to_float(-0.750),to_float(0.125),to_float(0.625),to_float(0.750),to_float(0.000),to_float(0.250),to_float(0.125),to_float(0.250),to_float(-0.750),to_float(0.250),to_float(0.875),to_float(0.375),to_float(-0.125),to_float(-0.375),to_float(0.625),to_float(-0.125)),
    (to_float(0.375),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(-0.125),to_float(0.625),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(-0.750),to_float(0.250),to_float(0.000),to_float(0.125),to_float(0.000)),
    (to_float(0.875),to_float(-0.875),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(-0.375),to_float(0.375),to_float(-0.875),to_float(-0.750),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(-0.625),to_float(0.875),to_float(-0.875)),
    (to_float(0.875),to_float(0.125),to_float(-0.375),to_float(0.625),to_float(-0.750),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.500),to_float(0.625),to_float(0.625),to_float(0.500),to_float(0.375),to_float(-0.375),to_float(0.875),to_float(-0.875)),
    (to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.125),to_float(-0.250),to_float(0.875),to_float(0.250),to_float(0.750),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(-0.375),to_float(0.500),to_float(0.875),to_float(0.625),to_float(-0.375),to_float(0.125),to_float(0.000),to_float(0.750),to_float(0.375)),
    (to_float(0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(0.750),to_float(0.000),to_float(-0.750),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.125)),
    (to_float(-0.125),to_float(-0.625),to_float(-0.625),to_float(0.375),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.250),to_float(0.125),to_float(0.750),to_float(-0.125),to_float(0.000),to_float(0.000)),
    (to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.375),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.875),to_float(0.875),to_float(0.750),to_float(0.875),to_float(0.500),to_float(0.000)),
    (to_float(-0.125),to_float(0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(-0.875)),
    (to_float(0.500),to_float(-0.125),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(-0.250),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.625),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.625),to_float(0.750),to_float(0.375),to_float(-0.875)),
    (to_float(0.625),to_float(-0.875),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.625),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.250),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(-0.375)),
    (to_float(-0.625),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(-0.500),to_float(-0.375),to_float(-0.375),to_float(-0.875),to_float(-0.625),to_float(0.125),to_float(0.375),to_float(-0.500),to_float(-0.750),to_float(0.250),to_float(0.000),to_float(0.875),to_float(-0.500),to_float(-0.250),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(-0.500),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(-0.375),to_float(-0.125),to_float(0.250),to_float(-0.875),to_float(-0.625),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.375),to_float(-0.625),to_float(-0.750),to_float(0.375)),
    (to_float(0.625),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.500),to_float(0.500),to_float(0.250),to_float(0.500),to_float(-0.500),to_float(0.625),to_float(0.000),to_float(-0.125),to_float(0.375),to_float(0.500),to_float(0.000),to_float(0.750),to_float(-0.125)),
    (to_float(0.250),to_float(-0.375),to_float(0.375),to_float(0.375),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(0.000),to_float(0.125),to_float(0.500),to_float(-0.250),to_float(0.125),to_float(-0.125),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(0.375),to_float(0.500),to_float(0.250)),
    (to_float(0.250),to_float(-0.250),to_float(0.500),to_float(0.625),to_float(0.000),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(-0.500),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.375),to_float(0.625),to_float(0.250),to_float(0.000),to_float(0.625),to_float(0.000),to_float(0.875),to_float(-0.125)),
    (to_float(-0.250),to_float(0.250),to_float(0.625),to_float(-0.500),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(-0.375),to_float(-0.500),to_float(0.625),to_float(0.500),to_float(0.125),to_float(0.125),to_float(0.250),to_float(-0.500)),
    (to_float(-0.375),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.250),to_float(0.000),to_float(0.375),to_float(0.125),to_float(0.375),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.500),to_float(-0.625)),
    (to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(0.250),to_float(0.625),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.875),to_float(0.250)),
    (to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.625),to_float(-0.625),to_float(-0.250),to_float(0.625),to_float(-0.875)),
    (to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(-0.250),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.375),to_float(-0.750),to_float(0.125),to_float(0.625),to_float(0.000)),
    (to_float(-0.125),to_float(-0.375),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(0.625),to_float(0.250),to_float(0.500),to_float(0.250),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(-0.625),to_float(-0.375),to_float(-0.125),to_float(0.250),to_float(-0.625),to_float(0.250),to_float(0.125)),
    (to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.625),to_float(0.750),to_float(0.125),to_float(0.625),to_float(0.250),to_float(-0.250),to_float(0.000),to_float(0.625),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(-0.250),to_float(0.500),to_float(0.125),to_float(0.250),to_float(0.250),to_float(0.750)),
    (to_float(-0.375),to_float(0.125),to_float(0.125),to_float(-0.750),to_float(0.375),to_float(0.000),to_float(0.875),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.125)),
    (to_float(-0.375),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.125),to_float(0.875),to_float(-0.250),to_float(0.500),to_float(0.125),to_float(0.375),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(0.500)),
    (to_float(-0.500),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.250),to_float(0.875),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(0.250),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.125)),
    (to_float(0.125),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.625),to_float(0.375),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(0.375),to_float(0.000),to_float(0.500),to_float(0.125),to_float(0.250),to_float(0.375)),
    (to_float(0.750),to_float(0.125),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.750),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.500),to_float(0.500)),
    (to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.750),to_float(-0.625),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.500),to_float(0.125),to_float(0.375),to_float(-0.625),to_float(0.375),to_float(0.500)),
    (to_float(-0.500),to_float(0.500),to_float(0.625),to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(-0.625),to_float(-0.375),to_float(-0.875),to_float(-0.500),to_float(-0.750),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(-0.500),to_float(0.375),to_float(0.500),to_float(0.125),to_float(0.750),to_float(-0.625)),
    (to_float(0.000),to_float(0.500),to_float(-0.500),to_float(0.750),to_float(-0.875),to_float(0.500),to_float(-0.500),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(-0.750),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.500)),
    (to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.625),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.750),to_float(-0.375),to_float(0.750),to_float(0.250),to_float(0.750),to_float(-0.125)),
    (to_float(0.875),to_float(-0.375),to_float(0.375),to_float(0.875),to_float(0.500),to_float(-0.375),to_float(0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.750),to_float(0.250),to_float(0.375),to_float(-0.375),to_float(-0.875)),
    (to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.875),to_float(0.375),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.625),to_float(0.250),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(-0.125),to_float(-0.875),to_float(0.375)),
    (to_float(0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.125),to_float(-0.125),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.125),to_float(0.875)),
    (to_float(0.625),to_float(-0.125),to_float(0.750),to_float(0.500),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(0.250),to_float(0.375),to_float(0.625),to_float(0.750),to_float(0.750),to_float(-0.625),to_float(0.375),to_float(0.750)),
    (to_float(0.125),to_float(0.875),to_float(0.375),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.875),to_float(0.500),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.125),to_float(-0.250),to_float(-0.750)),
    (to_float(0.125),to_float(-0.375),to_float(0.000),to_float(0.125),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(-0.125),to_float(-0.250),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(-0.500),to_float(-0.250),to_float(-0.375)),
    (to_float(0.625),to_float(0.875),to_float(0.000),to_float(0.250),to_float(0.500),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(-0.500),to_float(0.375),to_float(0.125),to_float(0.500),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.500),to_float(-0.500),to_float(0.500),to_float(-0.500),to_float(0.000)),
    (to_float(0.625),to_float(0.000),to_float(0.000),to_float(-0.625),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.750),to_float(-0.500),to_float(-0.250),to_float(-0.125),to_float(-0.500),to_float(-0.250),to_float(0.375),to_float(0.375),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(-0.125),to_float(0.125)),
    (to_float(-0.125),to_float(0.875),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(-0.375),to_float(-0.625),to_float(0.375),to_float(0.500)),
    (to_float(0.500),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(0.500),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.750),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(0.500),to_float(0.375)),
    (to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(0.875),to_float(-0.250),to_float(0.500),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(0.125),to_float(0.125),to_float(0.500),to_float(-0.500),to_float(0.500),to_float(0.250),to_float(-0.250),to_float(0.500),to_float(0.375)),
    (to_float(0.000),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(0.750),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.500),to_float(-0.125),to_float(0.500),to_float(0.625),to_float(0.375),to_float(0.500),to_float(0.375),to_float(0.125),to_float(0.750),to_float(0.250)),
    (to_float(-0.375),to_float(-0.375),to_float(0.625),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.875),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(0.875),to_float(0.125)),
    (to_float(0.000),to_float(-0.500),to_float(0.500),to_float(-0.375),to_float(0.000),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(0.250),to_float(0.125),to_float(0.375),to_float(-0.750),to_float(-0.125),to_float(0.500),to_float(-0.250)),
    (to_float(-0.125),to_float(0.000),to_float(-0.375),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(0.500),to_float(0.750),to_float(0.375),to_float(-0.375),to_float(-0.125),to_float(0.625),to_float(0.375),to_float(0.000),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.000),to_float(0.125)),
    (to_float(0.125),to_float(-0.250),to_float(0.375),to_float(-0.625),to_float(0.250),to_float(0.250),to_float(0.500),to_float(0.500),to_float(0.750),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.500),to_float(0.250),to_float(0.000),to_float(0.250),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.125)),
    (to_float(0.125),to_float(0.125),to_float(0.500),to_float(-0.875),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(0.875),to_float(0.375)),
    (to_float(-0.125),to_float(-0.625),to_float(0.000),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.625),to_float(0.375),to_float(0.375),to_float(-0.250),to_float(-0.500),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.875),to_float(0.750)),
    (to_float(-0.125),to_float(0.500),to_float(-0.375),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(0.625),to_float(0.375),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.750),to_float(0.000)),
    (to_float(-0.375),to_float(0.375),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(-0.625),to_float(-0.250),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(0.250),to_float(0.500)),
    (to_float(0.500),to_float(-0.500),to_float(-0.625),to_float(-0.875),to_float(-0.250),to_float(-0.250),to_float(0.000),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(0.000),to_float(0.500),to_float(0.875),to_float(0.250),to_float(0.125),to_float(0.250),to_float(0.750),to_float(-0.125)),
    (to_float(0.125),to_float(-0.125),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(0.750),to_float(0.000),to_float(-0.500),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(-0.250),to_float(0.250),to_float(-0.125)),
    (to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.625),to_float(-0.500),to_float(0.250),to_float(-0.625),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(0.500)),
    (to_float(0.000),to_float(-0.250),to_float(-0.500),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(0.875),to_float(0.375),to_float(0.375),to_float(-0.750),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.875),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.500),to_float(-0.125)),
    (to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(-0.750),to_float(0.375),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(-0.375),to_float(-0.500),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(-0.500)),
    (to_float(0.875),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(-0.625),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.250),to_float(0.250),to_float(-0.250),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(0.625),to_float(0.625),to_float(0.125),to_float(-0.250)),
    (to_float(0.875),to_float(-0.500),to_float(0.500),to_float(-0.875),to_float(0.625),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.125),to_float(0.375),to_float(0.125),to_float(-0.375),to_float(-0.625),to_float(-0.625)),
    (to_float(0.875),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.875),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.000),to_float(0.375),to_float(0.375),to_float(-0.250),to_float(-0.250),to_float(0.750),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.875),to_float(-0.625),to_float(0.125),to_float(0.000)),
    (to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.375),to_float(-0.125),to_float(0.875),to_float(0.000),to_float(0.125),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.500),to_float(-0.250),to_float(0.750),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(-0.500),to_float(-0.125),to_float(0.875),to_float(-0.125),to_float(0.875)),
    (to_float(-0.125),to_float(0.750),to_float(0.625),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(0.375),to_float(-0.500),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.750),to_float(-0.500)),
    (to_float(-0.250),to_float(0.250),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(-0.375),to_float(-0.375),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(-0.750)),
    (to_float(-0.500),to_float(0.625),to_float(0.625),to_float(-0.625),to_float(0.250),to_float(0.250),to_float(-0.875),to_float(0.625),to_float(0.750),to_float(0.125),to_float(0.875),to_float(-0.500),to_float(-0.250),to_float(0.875),to_float(0.250),to_float(-0.750),to_float(0.625),to_float(-0.750),to_float(0.250),to_float(-0.875)),
    (to_float(0.625),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(0.500),to_float(0.750),to_float(0.625),to_float(-0.750),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.750),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.000)),
    (to_float(0.000),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(-0.375),to_float(0.500),to_float(-0.375),to_float(0.500),to_float(0.250),to_float(0.875),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(-0.250),to_float(-0.125),to_float(0.375),to_float(-0.500)),
    (to_float(0.375),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(-0.500),to_float(0.250),to_float(0.000),to_float(0.500),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(0.750),to_float(0.000),to_float(0.250),to_float(-0.250)),
    (to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(0.000),to_float(0.500),to_float(0.750),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(0.375),to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(-0.750),to_float(0.750),to_float(-0.375)),
    (to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(0.500),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(-0.375),to_float(0.625),to_float(0.000),to_float(0.500),to_float(0.250),to_float(0.250),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(0.125)),
    (to_float(0.375),to_float(-0.250),to_float(0.000),to_float(0.625),to_float(-0.500),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(-0.250),to_float(0.500),to_float(0.625),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(0.000),to_float(-0.750),to_float(0.125),to_float(0.125),to_float(0.750),to_float(-0.250)),
    (to_float(-0.875),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(0.375),to_float(0.000),to_float(-0.625),to_float(0.500),to_float(0.250),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(0.625),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.000),to_float(0.375),to_float(-0.375)),
    (to_float(-0.625),to_float(-0.125),to_float(0.625),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.750),to_float(0.250)),
    (to_float(-0.875),to_float(0.000),to_float(-0.500),to_float(-0.875),to_float(0.375),to_float(-0.250),to_float(-0.500),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.375),to_float(-0.250),to_float(-0.875),to_float(-0.125),to_float(0.250),to_float(-0.375)),
    (to_float(0.125),to_float(-0.250),to_float(0.000),to_float(-0.750),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(0.625),to_float(0.000),to_float(0.875),to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.500),to_float(-0.250)),
    (to_float(0.875),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.250),to_float(0.125),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(0.750),to_float(0.250)),
    (to_float(-0.125),to_float(0.250),to_float(-0.125),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(0.250),to_float(-0.625),to_float(0.750),to_float(0.250),to_float(0.625),to_float(-0.375),to_float(0.625),to_float(0.125),to_float(0.875),to_float(-0.625)),
    (to_float(0.125),to_float(-0.375),to_float(-0.500),to_float(-0.875),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.625),to_float(0.125),to_float(0.250),to_float(0.125),to_float(0.875),to_float(-0.750)),
    (to_float(0.125),to_float(0.500),to_float(0.250),to_float(-0.875),to_float(0.750),to_float(-0.625),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(0.000),to_float(0.000),to_float(-0.625),to_float(-0.250),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.375),to_float(0.875)),
    (to_float(0.500),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(0.500),to_float(-0.625),to_float(-0.875),to_float(-0.250),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(0.250),to_float(0.625)),
    (to_float(0.250),to_float(0.750),to_float(-0.500),to_float(-0.750),to_float(0.000),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.375),to_float(0.375),to_float(-0.500),to_float(0.625),to_float(0.125),to_float(-0.250),to_float(-0.125)),
    (to_float(-0.500),to_float(-0.500),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(-0.500),to_float(-0.125),to_float(0.500),to_float(-0.625),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.250),to_float(0.875),to_float(-0.250)),
    (to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.625),to_float(0.500),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(-0.625),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(0.250),to_float(0.875),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.500),to_float(-0.375)),
    (to_float(0.500),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(0.750),to_float(0.500),to_float(0.875),to_float(-0.250),to_float(-0.625),to_float(0.875),to_float(-0.500),to_float(0.250),to_float(0.750),to_float(0.125),to_float(0.750)),
    (to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(0.125),to_float(-0.125),to_float(-0.875),to_float(0.500),to_float(0.500),to_float(0.875),to_float(0.375),to_float(-0.500),to_float(-0.875),to_float(-0.625),to_float(-0.125)),
    (to_float(0.875),to_float(-0.750),to_float(-0.250),to_float(-0.375),to_float(-0.375),to_float(0.750),to_float(0.875),to_float(-0.625),to_float(-0.875),to_float(-0.375),to_float(0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.750),to_float(-0.750),to_float(-0.625),to_float(-0.250),to_float(-0.875),to_float(0.375)),
    (to_float(0.125),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(-0.375),to_float(0.375),to_float(0.500),to_float(-0.375),to_float(-0.250),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(0.625),to_float(0.875),to_float(-0.750),to_float(0.250),to_float(0.000)),
    (to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(-0.250),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.500)),
    (to_float(-0.250),to_float(-0.875),to_float(0.375),to_float(0.750),to_float(0.875),to_float(0.375),to_float(0.625),to_float(0.875),to_float(0.375),to_float(0.625),to_float(0.375),to_float(-0.875),to_float(0.125),to_float(0.500),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.500),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(-0.500),to_float(0.625),to_float(0.750),to_float(-0.875),to_float(-0.375),to_float(0.750),to_float(0.875),to_float(0.250),to_float(-0.625),to_float(0.000),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.875),to_float(-0.250)),
    (to_float(0.875),to_float(0.250),to_float(0.250),to_float(0.750),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(0.375),to_float(0.875),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(-0.500),to_float(0.250),to_float(-0.625)),
    (to_float(-0.500),to_float(0.625),to_float(0.875),to_float(0.625),to_float(-0.250),to_float(0.750),to_float(-0.125),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(-0.750),to_float(-0.250),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(0.250)),
    (to_float(0.250),to_float(0.750),to_float(0.375),to_float(0.250),to_float(0.375),to_float(0.500),to_float(-0.375),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(0.750),to_float(-0.875),to_float(0.125),to_float(0.750),to_float(-0.375),to_float(-0.875),to_float(-0.625),to_float(0.500),to_float(0.750),to_float(-0.500)),
    (to_float(0.375),to_float(0.250),to_float(-0.500),to_float(0.000),to_float(-0.250),to_float(0.250),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(-0.375),to_float(0.000),to_float(0.500),to_float(0.125)),
    (to_float(0.375),to_float(-0.750),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(-0.250),to_float(0.375),to_float(0.000),to_float(0.250),to_float(0.500),to_float(0.125),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(-0.125),to_float(0.375),to_float(0.375)),
    (to_float(0.625),to_float(-0.250),to_float(0.125),to_float(0.625),to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(0.000),to_float(-0.375),to_float(0.500),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(0.375)),
    (to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.375),to_float(-0.625),to_float(-0.250),to_float(0.375),to_float(0.125),to_float(0.125),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(0.500),to_float(-0.500)),
    (to_float(0.250),to_float(-0.125),to_float(-0.750),to_float(0.125),to_float(-0.750),to_float(0.250),to_float(-0.250),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(-0.250),to_float(0.250),to_float(0.750),to_float(-0.875),to_float(-0.125),to_float(-0.125),to_float(0.375),to_float(0.750)),
    (to_float(-0.250),to_float(-0.500),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.625),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(0.250),to_float(0.750),to_float(-0.875),to_float(0.000),to_float(0.625),to_float(-0.500),to_float(0.500)),
    (to_float(-0.875),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.125),to_float(-0.500),to_float(-0.250),to_float(-0.750),to_float(-0.375),to_float(0.500),to_float(-0.750),to_float(-0.875),to_float(-0.375),to_float(0.000),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.500),to_float(0.375),to_float(-0.500),to_float(-0.125),to_float(0.625),to_float(-0.375),to_float(0.125),to_float(0.000),to_float(-0.250),to_float(-0.625),to_float(0.500),to_float(0.500),to_float(-0.375),to_float(0.125),to_float(-0.500),to_float(-0.875),to_float(-0.750),to_float(-0.125),to_float(0.125)),
    (to_float(-0.250),to_float(-0.625),to_float(-0.375),to_float(0.000),to_float(0.625),to_float(-0.625),to_float(-0.750),to_float(0.375),to_float(0.125),to_float(0.125),to_float(0.500),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(0.500),to_float(0.000),to_float(-0.500),to_float(0.000)),
    (to_float(-0.375),to_float(0.125),to_float(-0.500),to_float(0.500),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(-0.625),to_float(0.500),to_float(0.000),to_float(0.500),to_float(-0.250),to_float(0.125),to_float(0.625),to_float(0.250),to_float(-0.250),to_float(0.250),to_float(0.250)),
    (to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.500),to_float(0.125)),
    (to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(0.375),to_float(0.500),to_float(0.625),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.875)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.500),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(-0.500),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.500),to_float(0.375),to_float(0.250),to_float(-0.375),to_float(0.250)),
    (to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(0.500),to_float(0.625),to_float(-0.875),to_float(-0.750),to_float(0.000),to_float(0.250),to_float(0.500),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.750),to_float(-0.250),to_float(0.250)),
    (to_float(-0.500),to_float(-0.125),to_float(-0.375),to_float(0.750),to_float(-0.250),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(-0.625),to_float(-0.250),to_float(-0.625),to_float(-0.125),to_float(-0.250),to_float(0.625),to_float(0.250),to_float(0.375),to_float(-0.125),to_float(-0.500),to_float(0.125)),
    (to_float(0.375),to_float(0.125),to_float(0.500),to_float(0.375),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(0.125),to_float(0.500),to_float(-0.500),to_float(0.500),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.250),to_float(-0.500),to_float(-0.500),to_float(-0.125)),
    (to_float(-0.375),to_float(0.500),to_float(0.625),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(-0.750),to_float(0.000),to_float(0.375),to_float(-0.750),to_float(-0.375),to_float(-0.500),to_float(-0.500),to_float(-0.250),to_float(-0.875),to_float(0.125)),
    (to_float(0.875),to_float(0.750),to_float(0.125),to_float(0.375),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.500),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(0.625),to_float(-0.875),to_float(-0.625)),
    (to_float(-0.625),to_float(-0.625),to_float(-0.625),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(0.250),to_float(0.750),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(0.250),to_float(0.875),to_float(-0.250),to_float(-0.500)),
    (to_float(0.625),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.625),to_float(-0.250),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(0.000),to_float(-0.750),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.000)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(-0.750),to_float(0.500),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.000)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.250),to_float(0.375),to_float(0.375),to_float(-0.375),to_float(-0.375),to_float(0.625),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(0.750),to_float(0.875),to_float(-0.375),to_float(0.250),to_float(0.000)),
    (to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.625),to_float(-0.875),to_float(0.125),to_float(0.750),to_float(-0.750),to_float(0.875),to_float(0.875)),
    (to_float(-0.500),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(0.125),to_float(0.500),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(-0.875),to_float(-0.750),to_float(-0.250),to_float(0.875),to_float(0.875)),
    (to_float(0.750),to_float(0.125),to_float(-0.750),to_float(0.500),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.500),to_float(-0.375),to_float(0.250),to_float(0.500),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.625),to_float(-0.875)),
    (to_float(-0.250),to_float(0.500),to_float(0.250),to_float(0.375),to_float(-0.500),to_float(-0.250),to_float(-0.250),to_float(0.375),to_float(0.250),to_float(0.625),to_float(0.000),to_float(0.125),to_float(0.625),to_float(0.250),to_float(0.125),to_float(-0.875),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(-0.250)),
    (to_float(0.625),to_float(0.000),to_float(0.500),to_float(0.000),to_float(-0.875),to_float(-0.125),to_float(0.750),to_float(0.375),to_float(-0.125),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.500),to_float(-0.500)),
    (to_float(-0.375),to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.500),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(-0.250),to_float(0.125),to_float(0.750),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(0.375),to_float(-0.875),to_float(-0.500),to_float(-0.375),to_float(-0.750),to_float(0.875)),
    (to_float(0.375),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(-0.625),to_float(0.375),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.375),to_float(-0.875),to_float(-0.500),to_float(0.125),to_float(0.125),to_float(0.625)),
    (to_float(0.750),to_float(0.125),to_float(-0.625),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(0.750),to_float(-0.125),to_float(-0.875),to_float(-0.125),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.375)),
    (to_float(0.250),to_float(0.500),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(-0.125),to_float(0.375),to_float(-0.375),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(-0.625),to_float(-0.875),to_float(0.125),to_float(-0.500),to_float(-0.625),to_float(0.250)),
    (to_float(0.375),to_float(0.000),to_float(-0.500),to_float(0.125),to_float(0.625),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.125),to_float(0.125),to_float(-0.750),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(0.625),to_float(-0.750),to_float(0.125),to_float(0.625)),
    (to_float(0.500),to_float(0.625),to_float(-0.500),to_float(-0.375),to_float(-0.750),to_float(0.500),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(0.750),to_float(0.250),to_float(0.125),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(-0.125),to_float(-0.375)),
    (to_float(-0.875),to_float(0.750),to_float(-0.250),to_float(0.125),to_float(0.250),to_float(0.250),to_float(0.000),to_float(0.125),to_float(-0.250),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(0.125),to_float(-0.500),to_float(-0.375),to_float(0.000),to_float(-0.250)),
    (to_float(-0.875),to_float(0.125),to_float(0.500),to_float(0.250),to_float(0.625),to_float(0.750),to_float(0.625),to_float(0.750),to_float(-0.500),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(0.250),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(0.750)),
    (to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.500),to_float(0.125),to_float(0.625),to_float(-0.125),to_float(-0.625),to_float(0.125),to_float(0.000),to_float(0.250),to_float(-0.500),to_float(-0.625),to_float(0.000),to_float(-0.125),to_float(-0.750),to_float(-0.250),to_float(-0.375)),
    (to_float(-0.750),to_float(-0.375),to_float(-0.250),to_float(0.625),to_float(-0.625),to_float(0.750),to_float(-0.375),to_float(0.250),to_float(-0.750),to_float(0.375),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(0.250),to_float(0.500),to_float(-0.375),to_float(-0.125),to_float(0.125),to_float(-0.500),to_float(0.125)),
    (to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(0.875),to_float(0.750),to_float(0.375),to_float(-0.875),to_float(0.125),to_float(-0.500),to_float(0.625),to_float(0.375),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.750),to_float(-0.625)),
    (to_float(-0.500),to_float(0.250),to_float(0.500),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.625),to_float(-0.125),to_float(-0.625),to_float(-0.250),to_float(0.500),to_float(-0.250),to_float(-0.875),to_float(-0.125)),
    (to_float(0.125),to_float(-0.375),to_float(0.375),to_float(0.750),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.875),to_float(0.125),to_float(0.000),to_float(0.375),to_float(-0.375),to_float(0.500),to_float(-0.125),to_float(-0.625)),
    (to_float(-0.500),to_float(0.125),to_float(-0.375),to_float(0.625),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.250),to_float(0.375),to_float(0.000),to_float(0.875),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(0.500)),
    (to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.875),to_float(0.625),to_float(-0.625),to_float(-0.875),to_float(0.125),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(-0.625),to_float(0.375)),
    (to_float(0.500),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(-0.125),to_float(0.750),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.750),to_float(0.250)),
    (to_float(0.250),to_float(0.250),to_float(-0.625),to_float(0.375),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(-0.750),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.500),to_float(-0.875),to_float(-0.125),to_float(0.250)),
    (to_float(0.375),to_float(0.875),to_float(0.250),to_float(0.875),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(0.750),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.625),to_float(-0.250),to_float(-0.500),to_float(0.875),to_float(0.875)),
    (to_float(0.500),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(-0.125),to_float(-0.250),to_float(-0.625),to_float(0.875),to_float(-0.250),to_float(0.875)),
    (to_float(0.875),to_float(-0.500),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(-0.875),to_float(0.000),to_float(-0.250),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(-0.750),to_float(0.500)),
    (to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(0.500),to_float(-0.500),to_float(-0.375),to_float(0.625),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(0.500),to_float(0.875),to_float(-0.375),to_float(0.375),to_float(0.000)),
    (to_float(-0.500),to_float(-0.500),to_float(0.250),to_float(0.875),to_float(0.625),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(-0.250)),
    (to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.750),to_float(-0.875),to_float(0.000),to_float(0.125),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.500),to_float(0.125),to_float(0.875)),
    (to_float(0.875),to_float(0.000),to_float(0.000),to_float(0.375),to_float(0.750),to_float(-0.375),to_float(-0.125),to_float(-0.625),to_float(-0.500),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(0.875)),
    (to_float(0.500),to_float(0.500),to_float(-0.875),to_float(0.250),to_float(0.500),to_float(-0.125),to_float(0.875),to_float(-0.375),to_float(0.375),to_float(0.375),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(-0.625),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(-0.625),to_float(-0.250),to_float(0.000)),
    (to_float(-0.250),to_float(0.375),to_float(-0.875),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(-0.500),to_float(0.375),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(-0.500),to_float(0.000),to_float(-0.500),to_float(0.000)),
    (to_float(0.125),to_float(0.375),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(-0.625),to_float(0.250),to_float(-0.375),to_float(-0.500),to_float(0.125),to_float(-0.750),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.375),to_float(0.125),to_float(0.625)),
    (to_float(0.625),to_float(0.000),to_float(0.000),to_float(0.375),to_float(0.250),to_float(-0.250),to_float(-0.500),to_float(0.625),to_float(0.250),to_float(0.125),to_float(-0.625),to_float(-0.625),to_float(0.250),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.375),to_float(-0.625),to_float(-0.500),to_float(-0.250)),
    (to_float(-0.250),to_float(0.375),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(-0.250),to_float(0.750),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.500),to_float(-0.375),to_float(-0.125),to_float(-0.875)),
    (to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(-0.500),to_float(0.125),to_float(-0.375),to_float(0.375),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(0.250),to_float(-0.500),to_float(0.250),to_float(-0.375),to_float(-0.500),to_float(0.250)),
    (to_float(0.375),to_float(-0.375),to_float(0.500),to_float(-0.250),to_float(0.125),to_float(0.625),to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.125),to_float(0.375),to_float(-0.375),to_float(-0.375),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.500)),
    (to_float(0.500),to_float(-0.375),to_float(0.625),to_float(0.500),to_float(0.250),to_float(0.375),to_float(0.500),to_float(0.250),to_float(-0.500),to_float(-0.250),to_float(0.875),to_float(0.750),to_float(-0.125),to_float(-0.875),to_float(-0.125),to_float(0.750),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.125)),
    (to_float(0.750),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(0.750),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(-0.500),to_float(0.125),to_float(-0.500),to_float(-0.250)),
    (to_float(0.250),to_float(-0.625),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.625),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(0.625),to_float(-0.125),to_float(0.875),to_float(0.250),to_float(-0.500),to_float(0.750),to_float(0.375),to_float(0.625),to_float(0.000),to_float(-0.375),to_float(0.125)),
    (to_float(-0.625),to_float(-0.625),to_float(0.375),to_float(0.500),to_float(0.625),to_float(0.750),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(-0.500),to_float(-0.375),to_float(0.500),to_float(0.500),to_float(0.875),to_float(-0.500),to_float(0.125),to_float(0.000),to_float(0.625),to_float(-0.375),to_float(-0.125)),
    (to_float(0.000),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(0.750),to_float(0.000),to_float(-0.375),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(-0.750),to_float(0.625),to_float(-0.875),to_float(-0.750),to_float(-0.625),to_float(0.500),to_float(-0.375),to_float(0.250),to_float(-0.500)),
    (to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.625),to_float(-0.375),to_float(0.250),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.125)),
    (to_float(-0.625),to_float(0.125),to_float(0.875),to_float(0.250),to_float(0.750),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.625),to_float(0.250),to_float(0.125)),
    (to_float(-0.625),to_float(0.000),to_float(-0.125),to_float(0.375),to_float(0.500),to_float(0.250),to_float(0.375),to_float(0.625),to_float(0.250),to_float(0.125),to_float(0.500),to_float(0.125),to_float(0.500),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(0.250),to_float(0.250),to_float(0.125),to_float(-0.375)),
    (to_float(-0.125),to_float(0.000),to_float(-0.750),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(-0.375),to_float(-0.250),to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(0.875),to_float(-0.750),to_float(0.500),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.250),to_float(0.125)),
    (to_float(-0.125),to_float(0.750),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(0.750),to_float(-0.250),to_float(0.625),to_float(0.125),to_float(0.625),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(-0.125)),
    (to_float(0.250),to_float(0.875),to_float(0.375),to_float(0.500),to_float(-0.375),to_float(-0.125),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(0.625),to_float(0.250),to_float(0.375),to_float(0.625),to_float(0.375),to_float(-0.750),to_float(0.250),to_float(0.125),to_float(0.375),to_float(-0.875),to_float(0.750)),
    (to_float(0.375),to_float(0.625),to_float(0.125),to_float(0.375),to_float(-0.750),to_float(-0.375),to_float(-0.875),to_float(-0.500),to_float(0.125),to_float(0.375),to_float(-0.125),to_float(-0.625),to_float(-0.875),to_float(-0.500),to_float(0.250),to_float(-0.875),to_float(0.375),to_float(0.125),to_float(0.125),to_float(0.625)),
    (to_float(0.000),to_float(0.500),to_float(-0.125),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(-0.125),to_float(-0.375),to_float(-0.125),to_float(0.875)),
    (to_float(0.875),to_float(0.750),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(-0.625),to_float(0.125),to_float(-0.500),to_float(0.750),to_float(0.125),to_float(-0.875),to_float(0.875)),
    (to_float(0.875),to_float(0.625),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(0.375),to_float(-0.750),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.625),to_float(0.250),to_float(-0.250),to_float(0.125),to_float(0.500),to_float(-0.875)),
    (to_float(0.000),to_float(0.500),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.750),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(-0.125)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.625),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(-0.875),to_float(-0.375),to_float(0.750)),
    (to_float(0.375),to_float(-0.875),to_float(-0.375),to_float(0.250),to_float(-0.500),to_float(0.750),to_float(-0.125),to_float(0.875),to_float(0.500),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(-0.750),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(0.625),to_float(-0.375),to_float(-0.875),to_float(0.250)),
    (to_float(-0.125),to_float(-0.500),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(0.000),to_float(-0.875),to_float(0.625)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(-0.875)),
    (to_float(0.875),to_float(0.000),to_float(0.500),to_float(0.750),to_float(0.625),to_float(-0.750),to_float(-0.500),to_float(0.500),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(-0.500),to_float(0.125)),
    (to_float(-0.250),to_float(0.125),to_float(0.000),to_float(0.375),to_float(0.875),to_float(-0.250),to_float(-0.625),to_float(0.625),to_float(0.500),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.625)),
    (to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(0.625),to_float(-0.250),to_float(-0.500),to_float(-0.125),to_float(-0.625),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(0.375),to_float(-0.875),to_float(0.000),to_float(-0.500),to_float(0.500),to_float(-0.250),to_float(-0.625),to_float(-0.875)),
    (to_float(-0.250),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.750),to_float(-0.125),to_float(0.000),to_float(-0.375),to_float(-0.375),to_float(-0.375),to_float(-0.375),to_float(-0.500),to_float(-0.875),to_float(-0.375),to_float(0.500),to_float(0.750),to_float(0.125),to_float(-0.125),to_float(0.875)),
    (to_float(0.125),to_float(0.125),to_float(-0.250),to_float(0.375),to_float(-0.250),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(0.375),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(-0.125),to_float(0.750),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(-0.375),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.625),to_float(-0.375),to_float(-0.750),to_float(-0.250),to_float(-0.250),to_float(0.500),to_float(0.250),to_float(0.125),to_float(-0.875),to_float(0.250),to_float(0.375),to_float(0.375),to_float(0.625),to_float(0.375),to_float(0.500)),
    (to_float(0.500),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.375),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(0.500),to_float(0.500),to_float(0.000),to_float(-0.875),to_float(0.375),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(0.125)),
    (to_float(0.250),to_float(0.250),to_float(0.375),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.375),to_float(-0.500),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(0.625),to_float(0.000),to_float(0.625),to_float(-0.250),to_float(0.000)),
    (to_float(0.500),to_float(0.000),to_float(0.375),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.500),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.125)),
    (to_float(0.875),to_float(-0.625),to_float(-0.625),to_float(-0.125),to_float(-0.500),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(-0.750),to_float(0.625),to_float(0.125),to_float(0.875),to_float(0.125),to_float(0.500),to_float(0.250),to_float(0.500),to_float(-0.250),to_float(0.250),to_float(-0.250),to_float(-0.125)),
    (to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(-0.375),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(-0.625),to_float(0.625),to_float(-0.750),to_float(0.375),to_float(0.250),to_float(0.875),to_float(-0.375),to_float(0.250),to_float(-0.500),to_float(0.500),to_float(0.375),to_float(0.000)),
    (to_float(-0.375),to_float(-0.500),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.250),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(0.375),to_float(0.375),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(0.500),to_float(-0.375)),
    (to_float(0.125),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.125),to_float(0.125),to_float(-0.625),to_float(-0.375),to_float(-0.250),to_float(0.750),to_float(0.625),to_float(-0.625),to_float(-0.250),to_float(0.500),to_float(0.125),to_float(-0.125),to_float(-0.250),to_float(0.250)),
    (to_float(0.000),to_float(0.625),to_float(-0.250),to_float(-0.125),to_float(-0.500),to_float(0.750),to_float(-0.250),to_float(0.500),to_float(-0.875),to_float(0.125),to_float(0.125),to_float(0.375),to_float(0.125),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(-0.250),to_float(0.500),to_float(0.250),to_float(-0.250)),
    (to_float(-0.250),to_float(0.000),to_float(-0.375),to_float(-0.250),to_float(0.000),to_float(0.000),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.500),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(0.500),to_float(0.250),to_float(0.250),to_float(0.000)),
    (to_float(0.000),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.750),to_float(-0.250),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.125)),
    (to_float(0.000),to_float(0.875),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(0.250),to_float(-0.500),to_float(-0.375),to_float(0.375),to_float(-0.500),to_float(0.750),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.375)),
    (to_float(0.250),to_float(0.500),to_float(0.125),to_float(0.000),to_float(-0.750),to_float(0.125),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.750),to_float(0.500),to_float(-0.250),to_float(0.375),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(0.250)),
    (to_float(0.875),to_float(0.875),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.500),to_float(0.500),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(0.250),to_float(-0.250),to_float(-0.125),to_float(-0.375),to_float(0.500),to_float(0.125)),
    (to_float(0.125),to_float(0.875),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(-0.875),to_float(0.875)),
    (to_float(-0.750),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(0.250),to_float(-0.625),to_float(0.500),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(-0.375),to_float(-0.500),to_float(-0.250),to_float(-0.375),to_float(0.625),to_float(-0.875),to_float(0.250)),
    (to_float(0.625),to_float(0.125),to_float(0.125),to_float(0.750),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(0.875),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(0.250),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.250)),
    (to_float(-0.375),to_float(-0.125),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(-0.250),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.625),to_float(-0.500),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(0.125)),
    (to_float(0.125),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(-0.875),to_float(-0.500),to_float(0.625),to_float(0.875)),
    (to_float(0.500),to_float(-0.125),to_float(0.875),to_float(-0.250),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.125),to_float(-0.500),to_float(0.750),to_float(-0.625),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(0.875)),
    (to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(0.875),to_float(-0.625),to_float(0.750),to_float(0.000)),
    (to_float(-0.375),to_float(0.250),to_float(0.875),to_float(0.375),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.625),to_float(0.875),to_float(-0.125),to_float(-0.875)),
    (to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(-0.875)),
    (to_float(0.125),to_float(-0.125),to_float(0.625),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(0.250),to_float(-0.625),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.125),to_float(0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(0.875),to_float(0.625),to_float(-0.875),to_float(0.500),to_float(0.750),to_float(0.625),to_float(0.000),to_float(0.625),to_float(0.375),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.375),to_float(0.125)),
    (to_float(0.750),to_float(-0.125),to_float(0.500),to_float(-0.250),to_float(-0.500),to_float(-0.875),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(0.375),to_float(0.375),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(-0.625),to_float(0.875)),
    (to_float(0.500),to_float(-0.375),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.500),to_float(-0.125),to_float(0.000),to_float(0.625),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.000),to_float(0.000),to_float(0.250),to_float(0.250)),
    (to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(-0.625),to_float(0.250),to_float(0.250),to_float(0.875),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(0.625),to_float(0.000),to_float(0.000)),
    (to_float(0.625),to_float(0.250),to_float(0.125),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(-0.125),to_float(-0.750),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.125),to_float(0.125),to_float(0.125),to_float(0.250)),
    (to_float(0.500),to_float(-0.250),to_float(0.375),to_float(0.500),to_float(-0.250),to_float(-0.875),to_float(-0.375),to_float(-0.375),to_float(-0.375),to_float(0.750),to_float(-0.250),to_float(0.250),to_float(-0.625),to_float(-0.750),to_float(-0.500),to_float(0.875),to_float(-0.125),to_float(0.500),to_float(0.500),to_float(-0.125)),
    (to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.500),to_float(0.375),to_float(-0.625),to_float(0.500),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.250),to_float(0.500),to_float(0.500),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(-0.125)),
    (to_float(0.625),to_float(0.000),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(0.750),to_float(0.500),to_float(0.250),to_float(0.000),to_float(0.375),to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(0.125)),
    (to_float(0.625),to_float(-0.875),to_float(0.250),to_float(-0.250),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(-0.500),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(-0.250),to_float(0.375),to_float(0.125),to_float(0.500),to_float(0.250),to_float(-0.125)),
    (to_float(-0.125),to_float(-0.375),to_float(-0.125),to_float(-0.375),to_float(-0.375),to_float(0.000),to_float(0.125),to_float(-0.500),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(0.500),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.625)),
    (to_float(0.500),to_float(0.375),to_float(-0.375),to_float(-0.125),to_float(0.125),to_float(0.750),to_float(0.125),to_float(0.500),to_float(0.125),to_float(0.250),to_float(0.000),to_float(0.625),to_float(0.250),to_float(0.750),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.250)),
    (to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.250),to_float(0.500),to_float(-0.125),to_float(0.625),to_float(-0.375),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.625)),
    (to_float(-0.125),to_float(0.000),to_float(0.375),to_float(0.125),to_float(-0.375),to_float(0.500),to_float(0.750),to_float(0.500),to_float(-0.750),to_float(0.250),to_float(0.500),to_float(0.250),to_float(0.375),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(0.500),to_float(-0.125),to_float(-0.500)),
    (to_float(0.500),to_float(0.000),to_float(0.125),to_float(-0.250),to_float(0.250),to_float(0.000),to_float(-0.750),to_float(0.625),to_float(-0.125),to_float(0.500),to_float(0.500),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(0.000)),
    (to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.500),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.750),to_float(0.000),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(-0.500),to_float(-0.625),to_float(-0.625),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(-0.125),to_float(0.125)),
    (to_float(0.250),to_float(0.625),to_float(0.000),to_float(-0.500),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.625),to_float(0.125),to_float(0.750),to_float(0.000),to_float(-0.875),to_float(0.375),to_float(-0.125),to_float(-0.125),to_float(0.625),to_float(0.250),to_float(0.250),to_float(0.375)),
    (to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(0.875),to_float(-0.625),to_float(0.375),to_float(0.500),to_float(0.250),to_float(0.375),to_float(-0.875),to_float(-0.500),to_float(-0.375),to_float(-0.125),to_float(0.125),to_float(0.625),to_float(0.750),to_float(0.500)),
    (to_float(0.000),to_float(-0.250),to_float(0.125),to_float(0.500),to_float(0.375),to_float(-0.625),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(-0.375)),
    (to_float(0.000),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.125),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.500),to_float(-0.625),to_float(0.125)),
    (to_float(-0.625),to_float(0.750),to_float(0.250),to_float(0.250),to_float(-0.750),to_float(0.750),to_float(-0.375),to_float(0.875),to_float(0.125),to_float(-0.375),to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.500),to_float(0.375),to_float(0.875),to_float(-0.375),to_float(-0.625),to_float(0.000)),
    (to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(-0.875),to_float(0.500),to_float(0.500),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.250),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(0.500)),
    (to_float(0.000),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.375),to_float(0.375),to_float(0.125),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(0.750),to_float(-0.875),to_float(0.375),to_float(0.000),to_float(-0.625),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.375)),
    (to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.875)),
    (to_float(-0.625),to_float(-0.875),to_float(-0.125),to_float(-0.750),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.375),to_float(0.625),to_float(0.625),to_float(-0.875),to_float(0.750)),
    (to_float(0.875),to_float(-0.750),to_float(-0.750),to_float(0.875),to_float(0.500),to_float(-0.250),to_float(0.875),to_float(-0.375),to_float(-0.375),to_float(-0.750),to_float(-0.125),to_float(-0.750),to_float(-0.875),to_float(-0.500),to_float(0.250),to_float(-0.125),to_float(0.875),to_float(-0.375),to_float(0.625),to_float(0.000)),
    (to_float(-0.125),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.875),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(0.750),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.500),to_float(0.875),to_float(0.125),to_float(-0.125),to_float(0.000)),
    (to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(-0.500),to_float(-0.875)),
    (to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.500),to_float(0.500),to_float(-0.125),to_float(-0.500),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.750),to_float(-0.125),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(-0.750),to_float(-0.750),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.500),to_float(0.500)),
    (to_float(0.125),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.500),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.375),to_float(0.000),to_float(0.125),to_float(0.875)),
    (to_float(0.750),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(0.500),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(-0.500),to_float(0.250),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(-0.375),to_float(0.250),to_float(-0.125),to_float(-0.125)),
    (to_float(0.125),to_float(-0.250),to_float(0.750),to_float(0.375),to_float(0.125),to_float(-0.875),to_float(0.500),to_float(-0.625),to_float(0.250),to_float(0.750),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.500),to_float(0.375),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(0.250)),
    (to_float(-0.250),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.250),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(-0.250),to_float(-0.375),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(0.500),to_float(-0.250),to_float(0.125)),
    (to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(-0.375),to_float(-0.625),to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(0.750),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(0.625),to_float(0.375),to_float(0.000),to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(0.625)),
    (to_float(0.125),to_float(-0.500),to_float(0.625),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(0.500),to_float(-0.375),to_float(-0.125),to_float(0.875),to_float(0.000),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(0.375),to_float(0.125),to_float(0.750),to_float(0.125),to_float(0.625)),
    (to_float(0.625),to_float(0.000),to_float(0.375),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(-0.500),to_float(0.000),to_float(0.125),to_float(0.625),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.750),to_float(0.125),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(0.250),to_float(-0.125)),
    (to_float(0.125),to_float(-0.500),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(0.125),to_float(-0.375),to_float(-0.750),to_float(0.125),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(-0.250)),
    (to_float(0.000),to_float(0.000),to_float(-0.375),to_float(-0.125),to_float(-0.375),to_float(0.500),to_float(0.000),to_float(0.500),to_float(-0.250),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.625),to_float(0.250),to_float(-0.250),to_float(0.375)),
    (to_float(0.875),to_float(0.875),to_float(-0.125),to_float(-0.125),to_float(-0.500),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(0.875),to_float(-0.500),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(0.250),to_float(0.125)),
    (to_float(0.250),to_float(0.375),to_float(-0.625),to_float(0.000),to_float(0.000),to_float(-0.375),to_float(-0.250),to_float(0.625),to_float(-0.625),to_float(0.500),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(-0.500)),
    (to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.375),to_float(0.500),to_float(-0.125),to_float(-0.125),to_float(0.625),to_float(-0.125),to_float(-0.250),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(-0.500),to_float(0.125)),
    (to_float(0.125),to_float(0.500),to_float(-0.250),to_float(0.250),to_float(-0.625),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.375),to_float(0.625),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(0.375),to_float(-0.125)),
    (to_float(0.000),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(-0.625),to_float(0.500),to_float(-0.375),to_float(-0.250),to_float(-0.250),to_float(0.625),to_float(0.750),to_float(-0.375),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(0.000)),
    (to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.875),to_float(0.000),to_float(-0.375),to_float(0.500),to_float(0.500),to_float(-0.625),to_float(0.375),to_float(0.000),to_float(-0.250),to_float(-0.125),to_float(0.625),to_float(0.625),to_float(0.375)),
    (to_float(0.125),to_float(0.250),to_float(0.125),to_float(-0.375),to_float(0.750),to_float(0.750),to_float(0.250),to_float(-0.125),to_float(-0.500),to_float(-0.750),to_float(0.625),to_float(0.000),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(0.000)),
    (to_float(-0.750),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(-0.750),to_float(0.500),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(-0.375),to_float(0.000),to_float(-0.875),to_float(0.500),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.125)),
    (to_float(-0.500),to_float(-0.125),to_float(0.750),to_float(0.000),to_float(-0.500),to_float(0.250),to_float(-0.500),to_float(0.750),to_float(-0.250),to_float(0.375),to_float(0.875),to_float(-0.500),to_float(-0.125),to_float(-0.375),to_float(-0.875),to_float(-0.625),to_float(0.125),to_float(-0.500),to_float(0.250),to_float(0.125)),
    (to_float(0.250),to_float(-0.250),to_float(0.500),to_float(0.250),to_float(-0.875),to_float(0.625),to_float(-0.500),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(-0.125),to_float(-0.875),to_float(-0.625),to_float(-0.250),to_float(0.750),to_float(0.625),to_float(0.000),to_float(-0.875),to_float(0.375),to_float(0.250)),
    (to_float(-0.875),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.375),to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(0.125),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.500),to_float(0.750)),
    (to_float(0.250),to_float(-0.500),to_float(-0.125),to_float(0.875),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(-0.625),to_float(-0.500),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(0.625),to_float(-0.750),to_float(-0.625),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.125)),
    (to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.625),to_float(0.375),to_float(0.750),to_float(0.000),to_float(0.875),to_float(-0.500),to_float(0.000)),
    (to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(-0.125),to_float(0.750),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.250)),
    (to_float(-0.250),to_float(0.875),to_float(-0.500),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(-0.500),to_float(-0.625),to_float(0.125),to_float(0.875),to_float(-0.125),to_float(0.375),to_float(0.000)),
    (to_float(-0.375),to_float(-0.875),to_float(0.125),to_float(0.750),to_float(0.375),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(-0.625),to_float(-0.125),to_float(-0.625),to_float(-0.750),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.000)),
    (to_float(0.625),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(-0.500),to_float(0.250),to_float(-0.875)),
    (to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.250),to_float(0.500),to_float(0.750),to_float(-0.750),to_float(-0.375),to_float(0.250),to_float(0.875),to_float(0.500),to_float(0.125),to_float(0.500),to_float(0.500),to_float(-0.375),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.125),to_float(0.750),to_float(0.125),to_float(0.875),to_float(-0.125),to_float(-0.750),to_float(-0.500),to_float(-0.750),to_float(-0.875),to_float(0.750),to_float(0.375),to_float(-0.875),to_float(-0.750),to_float(0.000),to_float(0.875),to_float(0.250),to_float(0.500),to_float(0.125),to_float(0.000)),
    (to_float(-0.375),to_float(-0.250),to_float(0.625),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.750),to_float(-0.625),to_float(0.000),to_float(-0.250),to_float(0.750),to_float(-0.875),to_float(-0.250),to_float(-0.375),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(-0.125),to_float(0.250)),
    (to_float(-0.375),to_float(0.750),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(-0.125),to_float(-0.625),to_float(-0.250),to_float(0.375),to_float(-0.375),to_float(-0.125),to_float(0.750),to_float(-0.125),to_float(-0.250),to_float(-0.250),to_float(0.875),to_float(0.250),to_float(0.250)),
    (to_float(-0.625),to_float(-0.125),to_float(0.750),to_float(-0.250),to_float(-0.375),to_float(-0.750),to_float(-0.250),to_float(0.125),to_float(-0.750),to_float(0.000),to_float(0.375),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.125)),
    (to_float(-0.625),to_float(0.000),to_float(0.750),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.750),to_float(-0.625),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(-0.125)),
    (to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(-0.875),to_float(-0.250),to_float(0.500),to_float(-0.125),to_float(0.625),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(-0.375),to_float(0.500)),
    (to_float(0.125),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(0.500),to_float(-0.875),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(-0.750),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000)),
    (to_float(-0.250),to_float(0.125),to_float(0.875),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(0.500),to_float(-0.125),to_float(0.625),to_float(0.250),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(0.625),to_float(0.500),to_float(0.375)),
    (to_float(0.500),to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(-0.375),to_float(-0.750),to_float(0.375),to_float(-0.625),to_float(0.375),to_float(0.875),to_float(0.125),to_float(0.250),to_float(0.500),to_float(0.625),to_float(0.500),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000)),
    (to_float(0.375),to_float(0.375),to_float(-0.375),to_float(-0.375),to_float(-0.250),to_float(-0.500),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.875),to_float(-0.500),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(-0.625),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(-0.125)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(0.375),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.500),to_float(-0.375)),
    (to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.250),to_float(0.125),to_float(0.500),to_float(0.375),to_float(-0.125),to_float(0.375),to_float(0.750),to_float(-0.500),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(0.500),to_float(-0.375),to_float(-0.375)),
    (to_float(0.625),to_float(0.625),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.750),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(0.375),to_float(-0.125),to_float(0.500),to_float(-0.750),to_float(0.250),to_float(-0.375),to_float(0.250),to_float(0.000),to_float(-0.125)),
    (to_float(0.125),to_float(0.250),to_float(0.375),to_float(0.000),to_float(-0.375),to_float(-0.125),to_float(-0.125),to_float(-0.500),to_float(-0.500),to_float(-0.250),to_float(0.875),to_float(-0.250),to_float(-0.750),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(0.875),to_float(0.125),to_float(0.250)),
    (to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.500),to_float(0.375),to_float(0.625),to_float(-0.125),to_float(-0.500),to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(-0.625),to_float(0.375),to_float(-0.250),to_float(0.125),to_float(-0.625),to_float(0.250),to_float(0.500),to_float(-0.375)),
    (to_float(0.000),to_float(0.250),to_float(0.500),to_float(0.250),to_float(-0.500),to_float(0.375),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(-0.500),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(-0.500),to_float(0.250),to_float(0.500),to_float(0.125),to_float(0.375),to_float(0.000),to_float(-0.750)),
    (to_float(-0.125),to_float(-0.375),to_float(0.250),to_float(0.375),to_float(0.500),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(0.625),to_float(-0.250),to_float(-0.750),to_float(-0.750),to_float(-0.375),to_float(0.125),to_float(-0.250),to_float(0.125),to_float(0.375),to_float(-0.125)),
    (to_float(-0.750),to_float(0.250),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(0.625),to_float(-0.250),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(0.375),to_float(-0.875),to_float(-0.125),to_float(0.500),to_float(0.375),to_float(0.000),to_float(0.625),to_float(0.500),to_float(-0.250),to_float(0.375)),
    (to_float(-0.500),to_float(0.500),to_float(-0.125),to_float(0.500),to_float(-0.125),to_float(0.875),to_float(0.250),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(-0.875),to_float(0.375),to_float(0.375),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(0.000),to_float(-0.125)),
    (to_float(-0.125),to_float(-0.125),to_float(0.625),to_float(0.500),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(0.500),to_float(-0.500),to_float(0.125),to_float(0.750),to_float(-0.875),to_float(0.375),to_float(0.250),to_float(0.625),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(-0.375)),
    (to_float(-0.875),to_float(-0.625),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.250),to_float(-0.250),to_float(-0.750),to_float(0.125),to_float(-0.500),to_float(-0.625),to_float(0.250),to_float(-0.750),to_float(0.625),to_float(-0.750),to_float(-0.250),to_float(0.125),to_float(-0.875)),
    (to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.500),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.625),to_float(0.500),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.500)),
    (to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.625),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.750)),
    (to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(0.500),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000)),
    (to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.625),to_float(-0.375),to_float(0.750),to_float(-0.500),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(0.000)),
    (to_float(-0.875),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(-0.875)),
    (to_float(0.625),to_float(0.000),to_float(-0.750),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(0.500),to_float(0.875),to_float(-0.500),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.500)),
    (to_float(0.250),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.500),to_float(-0.500),to_float(-0.500),to_float(-0.875),to_float(0.250),to_float(0.625),to_float(0.125),to_float(0.750),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(0.000),to_float(0.250)),
    (to_float(-0.500),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(-0.250),to_float(0.375),to_float(0.625),to_float(0.375),to_float(0.250),to_float(0.125),to_float(0.375),to_float(0.000)),
    (to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(-0.625),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(-0.750),to_float(0.500),to_float(0.000),to_float(-0.250),to_float(0.375),to_float(0.625),to_float(-0.375),to_float(0.250),to_float(0.750),to_float(0.375),to_float(-0.375)),
    (to_float(-0.375),to_float(-0.375),to_float(0.625),to_float(-0.250),to_float(0.750),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.250)),
    (to_float(0.250),to_float(-0.250),to_float(0.125),to_float(0.500),to_float(-0.125),to_float(-0.500),to_float(0.625),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(0.125),to_float(0.125),to_float(-0.375),to_float(0.625),to_float(0.125),to_float(0.250)),
    (to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(-0.250),to_float(-0.500),to_float(-0.750),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.750)),
    (to_float(-0.125),to_float(-0.750),to_float(0.500),to_float(-0.125),to_float(0.125),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.875),to_float(0.750),to_float(0.375),to_float(0.375),to_float(0.000),to_float(-0.500),to_float(-0.750),to_float(0.500),to_float(0.500),to_float(0.000)),
    (to_float(0.625),to_float(0.375),to_float(0.625),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(0.625),to_float(0.500),to_float(0.000),to_float(0.000),to_float(0.500),to_float(-0.250),to_float(0.125)),
    (to_float(-0.375),to_float(0.875),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(-0.875),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.500),to_float(-0.875),to_float(0.250),to_float(0.375),to_float(0.625),to_float(-0.125),to_float(0.125),to_float(0.625),to_float(-0.125),to_float(-0.625),to_float(0.000)),
    (to_float(0.500),to_float(0.250),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(-0.875),to_float(-0.625),to_float(0.250),to_float(0.000),to_float(0.875),to_float(-0.250),to_float(-0.625),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(-0.625),to_float(0.250),to_float(0.125),to_float(-0.750)),
    (to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.625),to_float(0.750),to_float(-0.500),to_float(0.125),to_float(-0.500),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(-0.500),to_float(-0.375),to_float(0.000)),
    (to_float(0.125),to_float(0.375),to_float(-0.500),to_float(-0.250),to_float(-0.500),to_float(0.000),to_float(-0.250),to_float(0.375),to_float(-0.500),to_float(0.125),to_float(0.250),to_float(0.125),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(0.375),to_float(0.000)),
    (to_float(0.375),to_float(0.125),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.625),to_float(-0.125),to_float(-0.250)),
    (to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(-0.375),to_float(-0.625),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(-0.250),to_float(-0.250)),
    (to_float(-0.250),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(-0.125),to_float(0.500),to_float(-0.125),to_float(0.000),to_float(-0.375),to_float(0.500),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(-0.500),to_float(0.250),to_float(0.500),to_float(0.375),to_float(-0.250),to_float(-0.375)),
    (to_float(-0.750),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(-0.250),to_float(-0.750),to_float(-0.250),to_float(-0.500),to_float(-0.250),to_float(-0.250),to_float(-0.625),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.500),to_float(-0.250),to_float(-0.500),to_float(0.125)),
    (to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(0.625),to_float(-0.250)),
    (to_float(-0.625),to_float(-0.125),to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(0.750),to_float(0.500),to_float(0.750),to_float(-0.500),to_float(-0.125),to_float(-0.625),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(0.375),to_float(-0.500),to_float(0.375),to_float(0.750),to_float(-0.500),to_float(0.000)),
    (to_float(0.625),to_float(0.125),to_float(0.375),to_float(-0.375),to_float(-0.750),to_float(0.500),to_float(0.875),to_float(0.125),to_float(0.375),to_float(-0.375),to_float(0.625),to_float(-0.250),to_float(-0.625),to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.250)),
    (to_float(0.250),to_float(-0.625),to_float(0.375),to_float(0.000),to_float(-0.875),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(-0.500),to_float(-0.375),to_float(0.000),to_float(0.625),to_float(0.125),to_float(0.125),to_float(0.750),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(-0.375),to_float(-0.500)),
    (to_float(0.125),to_float(0.875),to_float(-0.625),to_float(0.000),to_float(0.375),to_float(0.375),to_float(-0.250),to_float(0.500),to_float(0.375),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(-0.125),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.375)),
    (to_float(-0.500),to_float(0.875),to_float(0.125),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.750),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.125)),
    (to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(0.750),to_float(0.000),to_float(0.625),to_float(-0.875)),
    (to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.750)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.375),to_float(-0.375),to_float(0.500),to_float(0.125),to_float(-0.375),to_float(0.375),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.375),to_float(0.875),to_float(-0.625),to_float(0.250),to_float(0.250)),
    (to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.625),to_float(0.250),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.750),to_float(-0.500),to_float(0.875),to_float(-0.625),to_float(-0.500),to_float(0.000),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(0.500),to_float(-0.875),to_float(-0.500),to_float(-0.250),to_float(-0.125)),
    (to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.625),to_float(0.375),to_float(0.875),to_float(0.750),to_float(0.125),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.125),to_float(0.625),to_float(0.000),to_float(-0.250),to_float(-0.375),to_float(0.875),to_float(-0.125),to_float(-0.125)),
    (to_float(0.125),to_float(-0.375),to_float(0.125),to_float(0.500),to_float(0.000),to_float(0.250),to_float(0.500),to_float(0.000),to_float(-0.125),to_float(-0.750),to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.500),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(-0.625)),
    (to_float(0.625),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(-0.875),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.125)),
    (to_float(-0.500),to_float(0.250),to_float(0.375),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(0.375),to_float(-0.500),to_float(0.250),to_float(-0.875),to_float(-0.500),to_float(-0.625),to_float(-0.375),to_float(0.750),to_float(-0.125),to_float(-0.500),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(0.125)),
    (to_float(0.125),to_float(-0.625),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.875),to_float(-0.500),to_float(-0.500),to_float(-0.375),to_float(-0.750),to_float(0.875),to_float(-0.375),to_float(-0.250),to_float(0.125),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.875),to_float(-0.125),to_float(0.375)),
    (to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.500),to_float(-0.375),to_float(-0.875),to_float(-0.375),to_float(0.625),to_float(-0.125),to_float(0.250),to_float(0.500),to_float(0.375),to_float(0.250),to_float(0.750),to_float(0.000),to_float(0.875)),
    (to_float(0.125),to_float(0.125),to_float(0.125),to_float(-0.375),to_float(0.000),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(-0.500),to_float(-0.625),to_float(-0.375),to_float(0.500),to_float(0.500),to_float(-0.625),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.375)),
    (to_float(-0.250),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.500),to_float(-0.500),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.000)),
    (to_float(0.250),to_float(0.875),to_float(-0.250),to_float(-0.500),to_float(-0.250),to_float(-0.875),to_float(0.625),to_float(-0.250),to_float(-0.500),to_float(0.000),to_float(-0.875),to_float(0.625),to_float(0.375),to_float(0.375),to_float(0.125),to_float(0.000),to_float(0.625),to_float(0.375),to_float(-0.250),to_float(-0.875)),
    (to_float(0.875),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(0.625),to_float(-0.625),to_float(-0.500),to_float(0.500),to_float(-0.875),to_float(-0.125),to_float(-0.625),to_float(0.000),to_float(-0.250),to_float(0.375),to_float(-0.500),to_float(-0.625),to_float(0.375),to_float(0.625),to_float(0.125),to_float(-0.250)),
    (to_float(0.000),to_float(0.125),to_float(-0.375),to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.250),to_float(0.375),to_float(-0.250),to_float(0.125),to_float(0.875),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(0.875),to_float(0.375),to_float(0.250)),
    (to_float(-0.500),to_float(0.500),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(-0.250)),
    (to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.500),to_float(0.250),to_float(0.500),to_float(0.375),to_float(-0.875),to_float(0.000),to_float(-0.250),to_float(0.750),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.000),to_float(-0.125)),
    (to_float(-0.375),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.500),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(0.375),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(0.125)),
    (to_float(-0.625),to_float(0.375),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.125),to_float(0.500),to_float(0.000),to_float(-0.375),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.125),to_float(-0.250)),
    (to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.500),to_float(-0.500),to_float(0.750),to_float(0.125),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.500),to_float(0.250),to_float(-0.375),to_float(-0.375)),
    (to_float(0.000),to_float(-0.125),to_float(-0.375),to_float(-0.625),to_float(-0.625),to_float(0.250),to_float(0.375),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(-0.500),to_float(0.000),to_float(-0.750),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(-0.500),to_float(0.375),to_float(0.250)),
    (to_float(-0.625),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(-0.875),to_float(0.375),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.500),to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(0.500),to_float(0.500),to_float(-0.125),to_float(-0.250),to_float(-0.125)),
    (to_float(-0.250),to_float(0.250),to_float(0.625),to_float(-0.500),to_float(-0.875),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(-0.750),to_float(-0.375),to_float(0.125),to_float(-0.500),to_float(-0.250),to_float(0.625),to_float(0.125)),
    (to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(-0.500),to_float(0.750),to_float(-0.125),to_float(0.375),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(0.000),to_float(-0.500),to_float(-0.500),to_float(0.375),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125)),
    (to_float(0.000),to_float(-0.875),to_float(-0.250),to_float(-0.375),to_float(0.375),to_float(0.000),to_float(-0.750),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(0.875),to_float(0.000),to_float(-0.250),to_float(-0.875),to_float(-0.625),to_float(-0.875),to_float(0.875)),
    (to_float(0.875),to_float(-0.750),to_float(-0.750),to_float(0.250),to_float(0.750),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.875)),
    (to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.125)),
    (to_float(0.250),to_float(-0.875),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.750),to_float(-0.250),to_float(0.375),to_float(0.625),to_float(-0.250),to_float(0.125),to_float(0.875),to_float(-0.375),to_float(0.000),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.000),to_float(0.625)),
    (to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.125),to_float(0.500),to_float(0.750),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.250),to_float(0.750),to_float(-0.250)),
    (to_float(0.250),to_float(-0.875),to_float(0.375),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(-0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(-0.125),to_float(0.000),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.375),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.625),to_float(-0.375),to_float(-0.625),to_float(-0.625),to_float(-0.250),to_float(0.250),to_float(-0.500)),
    (to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.375),to_float(-0.500),to_float(-0.375),to_float(0.875),to_float(-0.625),to_float(-0.375)),
    (to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(0.375),to_float(0.625),to_float(0.500),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(0.375),to_float(0.125),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(0.000)),
    (to_float(-0.250),to_float(0.000),to_float(0.500),to_float(-0.375),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(-0.625),to_float(0.750),to_float(-0.250),to_float(-0.250),to_float(0.000)),
    (to_float(0.125),to_float(-0.500),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.125),to_float(-0.875),to_float(-0.625),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(-0.250),to_float(0.250)),
    (to_float(-0.125),to_float(-0.625),to_float(0.125),to_float(-0.250),to_float(0.250),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.625),to_float(-0.500),to_float(0.500),to_float(0.875)),
    (to_float(0.000),to_float(0.375),to_float(0.750),to_float(0.500),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.500),to_float(-0.750),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(0.875)),
    (to_float(0.125),to_float(0.500),to_float(-0.375),to_float(0.250),to_float(-0.625),to_float(-0.250),to_float(0.375),to_float(0.125),to_float(0.125),to_float(-0.875),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(0.250),to_float(0.375),to_float(0.750),to_float(-0.250),to_float(-0.875)),
    (to_float(-0.250),to_float(0.625),to_float(0.000),to_float(-0.375),to_float(-0.125),to_float(-0.375),to_float(0.500),to_float(0.125),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(-0.375),to_float(-0.375),to_float(0.625),to_float(0.750),to_float(-0.750),to_float(0.000),to_float(0.750),to_float(-0.250)),
    (to_float(0.875),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(0.375),to_float(-0.250),to_float(-0.250),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.625),to_float(-0.125),to_float(-0.125),to_float(0.375),to_float(-0.500),to_float(0.750),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(0.000)),
    (to_float(0.500),to_float(-0.125),to_float(0.625),to_float(0.250),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(0.625),to_float(0.250),to_float(-0.250),to_float(-0.500),to_float(0.875),to_float(0.250),to_float(0.000)),
    (to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.250),to_float(0.125),to_float(-0.375),to_float(0.000),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(0.500),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.500),to_float(-0.250),to_float(-0.250)),
    (to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(0.000),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(-0.250),to_float(-0.625),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(-0.500),to_float(0.000)),
    (to_float(0.000),to_float(0.250),to_float(0.375),to_float(0.000),to_float(0.250),to_float(0.125),to_float(0.250),to_float(-0.375),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(-0.500),to_float(0.000),to_float(0.250),to_float(0.250),to_float(0.375),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(-0.125)),
    (to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.125),to_float(0.750),to_float(0.125),to_float(0.375),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(-0.500),to_float(0.125),to_float(-0.125),to_float(-0.125)),
    (to_float(-0.625),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(-0.500),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(0.250),to_float(0.625),to_float(0.125)),
    (to_float(0.625),to_float(-0.375),to_float(-0.375),to_float(0.000),to_float(-0.750),to_float(-0.375),to_float(-0.375),to_float(-0.500),to_float(0.250),to_float(-0.375),to_float(-0.500),to_float(-0.125),to_float(0.250),to_float(-0.625),to_float(-0.250),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(-0.250),to_float(-0.250)),
    (to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(-0.875),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.375),to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(0.125),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(0.375)),
    (to_float(-0.500),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(-0.625),to_float(-0.250),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(-0.500),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(-0.375),to_float(0.250),to_float(0.250)),
    (to_float(0.750),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(0.750),to_float(0.125),to_float(0.625),to_float(-0.375),to_float(-0.500),to_float(-0.875),to_float(-0.500),to_float(0.750),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(0.000)),
    (to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(-0.625),to_float(-0.250),to_float(0.875),to_float(-0.500),to_float(0.375),to_float(0.125),to_float(-0.875),to_float(-0.125)),
    (to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.000),to_float(0.375),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(-0.625)),
    (to_float(0.000),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(-0.875),to_float(0.875)),
    (to_float(0.875),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.125),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(0.875)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.125)),
    (to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.250),to_float(0.375),to_float(-0.750),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.750),to_float(-0.875),to_float(-0.500),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(-0.875)),
    (to_float(-0.250),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(0.750),to_float(-0.750),to_float(0.375),to_float(-0.875),to_float(0.375),to_float(-0.125),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(0.750),to_float(0.125),to_float(-0.125),to_float(-0.500),to_float(-0.125),to_float(0.000),to_float(0.625),to_float(-0.375)),
    (to_float(-0.625),to_float(-0.375),to_float(0.000),to_float(-0.750),to_float(-0.250),to_float(0.625),to_float(0.750),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.000),to_float(-0.875),to_float(-0.125),to_float(0.625),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.125),to_float(0.875)),
    (to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.250),to_float(0.000),to_float(0.375),to_float(-0.250),to_float(-0.750),to_float(0.875),to_float(0.500),to_float(0.375),to_float(0.375),to_float(0.125),to_float(0.875),to_float(0.750),to_float(-0.625),to_float(0.250),to_float(-0.625),to_float(-0.625),to_float(0.125)),
    (to_float(0.125),to_float(0.125),to_float(0.625),to_float(-0.750),to_float(0.125),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(-0.625),to_float(-0.625),to_float(0.000),to_float(-0.125),to_float(0.875),to_float(0.000),to_float(-0.125),to_float(0.500),to_float(0.500),to_float(0.250),to_float(-0.250)),
    (to_float(-0.250),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.625),to_float(0.500),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(-0.500),to_float(0.375),to_float(0.750),to_float(0.500),to_float(0.250),to_float(0.125),to_float(-0.375),to_float(0.000),to_float(0.500)),
    (to_float(0.250),to_float(0.375),to_float(0.125),to_float(0.375),to_float(-0.375),to_float(0.500),to_float(0.125),to_float(-0.625),to_float(0.375),to_float(-0.500),to_float(-0.875),to_float(0.125),to_float(-0.250),to_float(0.250),to_float(-0.375),to_float(0.375),to_float(0.250),to_float(0.500),to_float(-0.500),to_float(0.375)),
    (to_float(0.625),to_float(0.750),to_float(0.250),to_float(0.500),to_float(0.375),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.750),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(-0.500),to_float(0.250),to_float(0.375)),
    (to_float(0.125),to_float(0.250),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(0.750),to_float(0.125),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(0.375),to_float(0.500),to_float(-0.375),to_float(-0.250),to_float(0.000),to_float(-0.625),to_float(-0.875)),
    (to_float(-0.375),to_float(0.750),to_float(0.500),to_float(-0.250),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.250),to_float(0.500),to_float(-0.125),to_float(-0.250),to_float(-0.500),to_float(-0.625),to_float(-0.375)),
    (to_float(0.000),to_float(-0.250),to_float(0.000),to_float(0.250),to_float(0.750),to_float(0.250),to_float(0.500),to_float(-0.125),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(-0.375),to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(-0.375),to_float(-0.500)),
    (to_float(-0.125),to_float(-0.125),to_float(0.375),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(-0.125),to_float(-0.750),to_float(0.250),to_float(0.000),to_float(-0.250),to_float(0.000),to_float(-0.750)),
    (to_float(0.250),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(-0.750),to_float(-0.875),to_float(0.625),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.375),to_float(0.000),to_float(0.125),to_float(0.500),to_float(0.125),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(-0.125)),
    (to_float(0.375),to_float(0.000),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(-0.250),to_float(0.250),to_float(-0.375),to_float(-0.500),to_float(0.000),to_float(0.250),to_float(0.125),to_float(-0.250)),
    (to_float(0.000),to_float(-0.500),to_float(-0.125),to_float(0.125),to_float(0.750),to_float(0.000),to_float(-0.125),to_float(0.625),to_float(0.625),to_float(0.000),to_float(-0.250),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(-0.500),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.750)),
    (to_float(0.375),to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(-0.375),to_float(0.625),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.375),to_float(-0.875),to_float(-0.500),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.500),to_float(0.000),to_float(0.250),to_float(-0.250),to_float(0.000)),
    (to_float(-0.125),to_float(-0.625),to_float(-0.250),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(-0.625),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.375),to_float(-0.500)),
    (to_float(0.125),to_float(-0.125),to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(-0.625),to_float(0.000),to_float(0.625),to_float(-0.375),to_float(-0.875),to_float(0.125),to_float(0.750),to_float(0.125),to_float(-0.375),to_float(-0.250),to_float(-0.375),to_float(-0.500),to_float(-0.250),to_float(-0.750)),
    (to_float(0.125),to_float(-0.750),to_float(0.500),to_float(-0.250),to_float(-0.625),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.625),to_float(-0.125),to_float(-0.875),to_float(-0.750),to_float(0.000),to_float(0.500),to_float(0.875),to_float(0.125),to_float(-0.500),to_float(0.000),to_float(-0.375),to_float(0.250)),
    (to_float(-0.250),to_float(-0.250),to_float(-0.250),to_float(0.625),to_float(0.875),to_float(0.750),to_float(0.625),to_float(-0.250),to_float(-0.250),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.375),to_float(-0.500),to_float(0.375),to_float(0.000),to_float(-0.625),to_float(-0.875),to_float(0.125)),
    (to_float(-0.250),to_float(0.000),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(0.625),to_float(-0.250),to_float(0.250),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.125),to_float(0.250),to_float(-0.250),to_float(0.250),to_float(0.375),to_float(-0.750),to_float(0.250)),
    (to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(-0.625),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(-0.125),to_float(-0.500),to_float(0.000),to_float(-0.375),to_float(-0.875),to_float(0.500),to_float(0.500),to_float(-0.250)),
    (to_float(0.250),to_float(-0.750),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.625),to_float(0.875),to_float(-0.500),to_float(-0.500),to_float(0.000),to_float(-0.750),to_float(0.625),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.125)),
    (to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(-0.500),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.000),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(0.875)),
    (to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.375),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(0.875),to_float(-0.500),to_float(0.125),to_float(0.125)),
    (to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(0.000),to_float(-0.375),to_float(0.875),to_float(0.750),to_float(-0.375),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(0.375)),
    (to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(0.000),to_float(0.625),to_float(-0.500),to_float(0.250),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(0.250),to_float(0.000)),
    (to_float(-0.625),to_float(-0.750),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.750),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.625),to_float(-0.375)),
    (to_float(0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.625),to_float(-0.625),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(0.500),to_float(-0.500),to_float(-0.625),to_float(0.750)),
    (to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(0.625),to_float(0.625),to_float(0.250),to_float(0.250),to_float(0.750),to_float(-0.500),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(0.500)),
    (to_float(-0.375),to_float(-0.375),to_float(-0.875),to_float(0.000),to_float(-0.625),to_float(0.625),to_float(0.875),to_float(-0.375),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(-0.500),to_float(-0.250),to_float(-0.125),to_float(-0.750),to_float(-0.500),to_float(0.250),to_float(0.625),to_float(0.250)),
    (to_float(-0.125),to_float(0.250),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(-0.125),to_float(0.000),to_float(0.500),to_float(-0.125),to_float(-0.625),to_float(0.375),to_float(0.125),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.250),to_float(-0.375),to_float(0.250)),
    (to_float(0.500),to_float(-0.125),to_float(0.250),to_float(0.625),to_float(0.500),to_float(0.500),to_float(0.125),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(-0.250),to_float(0.625),to_float(-0.500),to_float(0.125),to_float(-0.625),to_float(0.500),to_float(0.375),to_float(0.375)),
    (to_float(0.250),to_float(0.750),to_float(0.250),to_float(0.375),to_float(-0.375),to_float(0.875),to_float(-0.625),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(-0.625)),
    (to_float(0.250),to_float(-0.250),to_float(0.000),to_float(-0.500),to_float(-0.250),to_float(0.625),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.625),to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(0.125)),
    (to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.375),to_float(0.375),to_float(0.625),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.500),to_float(0.250),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(0.625)),
    (to_float(0.000),to_float(-0.250),to_float(0.625),to_float(-0.125),to_float(-0.250),to_float(0.375),to_float(0.250),to_float(-0.375),to_float(0.500),to_float(0.625),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(0.000),to_float(0.125),to_float(-0.250),to_float(-0.500),to_float(-0.125)),
    (to_float(0.125),to_float(0.000),to_float(0.500),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.375)),
    (to_float(0.125),to_float(0.875),to_float(-0.500),to_float(0.000),to_float(-0.500),to_float(0.125),to_float(0.000),to_float(-0.500),to_float(0.750),to_float(-0.375),to_float(0.250),to_float(-0.125),to_float(-0.375),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(-0.125)),
    (to_float(0.250),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(0.875),to_float(-0.250),to_float(-0.625),to_float(-0.500),to_float(-0.250),to_float(-0.125),to_float(-0.750),to_float(-0.250),to_float(-0.500),to_float(-0.625),to_float(-0.125),to_float(-0.750)),
    (to_float(0.000),to_float(-0.125),to_float(0.500),to_float(0.125),to_float(-0.500),to_float(-0.250),to_float(-0.125),to_float(-0.500),to_float(0.250),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.500),to_float(-0.500),to_float(0.000),to_float(-0.625)),
    (to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(-0.375),to_float(-0.250),to_float(0.500),to_float(-0.375)),
    (to_float(0.375),to_float(0.875),to_float(-0.625),to_float(0.125),to_float(0.500),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(-0.500),to_float(-0.125),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(-0.375),to_float(0.000)),
    (to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(0.250),to_float(-0.625),to_float(0.250),to_float(-0.500),to_float(0.250),to_float(-0.250),to_float(0.000),to_float(-0.500),to_float(-0.125),to_float(-0.250),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.000),to_float(0.375),to_float(-0.625)),
    (to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(0.250),to_float(0.250),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(-0.500),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.625),to_float(-0.250),to_float(-0.625)),
    (to_float(0.250),to_float(-0.625),to_float(-0.125),to_float(0.250),to_float(-0.875),to_float(0.250),to_float(0.125),to_float(0.250),to_float(-0.500),to_float(-0.750),to_float(-0.750),to_float(0.000),to_float(-0.500),to_float(-0.500),to_float(-0.250),to_float(-0.625),to_float(0.125),to_float(-0.625),to_float(0.125),to_float(-0.750)),
    (to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(-0.250),to_float(0.250),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(-0.500),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(-0.625),to_float(-0.125),to_float(0.875),to_float(0.375),to_float(0.000)),
    (to_float(0.625),to_float(-0.625),to_float(0.125),to_float(0.000),to_float(-0.375),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.375),to_float(-0.125),to_float(-0.875),to_float(0.625),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.375),to_float(-0.500),to_float(0.875)),
    (to_float(0.875),to_float(-0.875),to_float(-0.625),to_float(-0.500),to_float(-0.375),to_float(-0.250),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(-0.875),to_float(-0.750)),
    (to_float(0.125),to_float(-0.250),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.750),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(-0.250),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.625)),
    (to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(0.625),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.875),to_float(0.000),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.250),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.875)),
    (to_float(-0.125),to_float(-0.625),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(-0.500),to_float(0.125),to_float(0.125),to_float(0.625),to_float(-0.125),to_float(0.000),to_float(0.125)),
    (to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(-0.125),to_float(-0.125),to_float(-0.500),to_float(0.750),to_float(0.625),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(0.750),to_float(-0.250),to_float(0.125),to_float(0.375)),
    (to_float(-0.125),to_float(-0.875),to_float(-0.500),to_float(0.500),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.500),to_float(-0.875),to_float(-0.500),to_float(-0.125),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(0.125),to_float(0.125)),
    (to_float(-0.625),to_float(-0.625),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(0.375),to_float(-0.625),to_float(0.125),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(-0.500),to_float(0.375)),
    (to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.375),to_float(-0.500),to_float(0.625),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.625),to_float(0.000),to_float(-0.500),to_float(0.875)),
    (to_float(0.250),to_float(-0.500),to_float(-0.375),to_float(-0.875),to_float(0.500),to_float(0.125),to_float(0.125),to_float(0.375),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(-0.375),to_float(0.625),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(-0.375),to_float(0.125),to_float(0.375)),
    (to_float(0.000),to_float(0.500),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(-0.125),to_float(0.250),to_float(-0.875),to_float(-0.250),to_float(-0.500),to_float(0.875),to_float(-0.125),to_float(0.250),to_float(0.250),to_float(-0.500),to_float(-0.250),to_float(0.375)),
    (to_float(-0.250),to_float(-0.875),to_float(0.625),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(-0.375),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(0.125),to_float(0.500),to_float(-0.625),to_float(0.125),to_float(-0.500),to_float(0.375),to_float(0.125),to_float(-0.750),to_float(0.125)),
    (to_float(0.000),to_float(-0.250),to_float(0.125),to_float(-0.625),to_float(0.250),to_float(-0.250),to_float(0.500),to_float(0.375),to_float(0.250),to_float(0.125),to_float(-0.625),to_float(-0.500),to_float(0.500),to_float(-0.125),to_float(0.375),to_float(0.250),to_float(0.375),to_float(-0.250),to_float(-0.375),to_float(0.250)),
    (to_float(-0.250),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(0.000),to_float(0.375),to_float(0.250),to_float(0.625),to_float(0.375),to_float(0.750),to_float(0.000),to_float(0.125),to_float(0.500),to_float(0.000),to_float(0.125),to_float(0.375),to_float(-0.750),to_float(-0.375),to_float(0.625)),
    (to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(0.500),to_float(-0.375),to_float(-0.125),to_float(0.000),to_float(0.875),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(-0.625),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(0.000),to_float(-0.500),to_float(-0.375),to_float(0.250)),
    (to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(-0.250),to_float(-0.250),to_float(0.500),to_float(0.250),to_float(-0.375),to_float(0.125),to_float(0.125),to_float(0.875)),
    (to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.750),to_float(-0.125),to_float(0.000),to_float(0.375),to_float(0.750),to_float(0.375),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(-0.750),to_float(-0.250)),
    (to_float(0.250),to_float(0.000),to_float(0.375),to_float(0.125),to_float(0.375),to_float(-0.375),to_float(0.250),to_float(-0.500),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(-0.125),to_float(-0.250),to_float(0.375)),
    (to_float(0.000),to_float(0.375),to_float(-0.125),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(0.375),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(-0.875),to_float(-0.250)),
    (to_float(0.250),to_float(-0.500),to_float(-0.125),to_float(-0.125),to_float(0.750),to_float(0.250),to_float(0.250),to_float(0.000),to_float(0.375),to_float(-0.625),to_float(0.625),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(-0.250),to_float(-0.125),to_float(-0.375),to_float(-0.625),to_float(0.000),to_float(-0.250)),
    (to_float(-0.125),to_float(0.125),to_float(0.625),to_float(-0.250),to_float(0.500),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.375),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(0.000),to_float(-0.250),to_float(0.250),to_float(0.125),to_float(0.125),to_float(-0.500),to_float(-0.750),to_float(-0.875)),
    (to_float(-0.125),to_float(-0.500),to_float(0.125),to_float(-0.125),to_float(-0.625),to_float(-0.125),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(-0.375),to_float(0.125),to_float(0.000),to_float(-0.500),to_float(-0.250),to_float(-0.750),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(0.000),to_float(-0.250)),
    (to_float(0.125),to_float(-0.375),to_float(0.375),to_float(0.250),to_float(-0.500),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(-0.500),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(-0.500),to_float(-0.250),to_float(-0.250)),
    (to_float(0.125),to_float(-0.250),to_float(-0.625),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(0.000),to_float(0.375),to_float(0.375),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(0.000),to_float(0.250),to_float(0.125),to_float(-0.375),to_float(-0.500),to_float(-0.250),to_float(0.000),to_float(-0.125)),
    (to_float(0.625),to_float(-0.375),to_float(0.500),to_float(-0.250),to_float(-0.875),to_float(-0.375),to_float(0.500),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(0.500),to_float(-0.250),to_float(0.625),to_float(0.000),to_float(0.000),to_float(-0.500),to_float(-0.250)),
    (to_float(-0.375),to_float(-0.125),to_float(-0.750),to_float(-0.625),to_float(-0.875),to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.750),to_float(0.125),to_float(-0.375),to_float(0.125),to_float(0.250),to_float(0.500),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(-0.625)),
    (to_float(0.375),to_float(-0.125),to_float(0.250),to_float(-0.625),to_float(-0.500),to_float(-0.750),to_float(-0.625),to_float(0.000),to_float(-0.375),to_float(-0.875),to_float(-0.750),to_float(-0.500),to_float(0.250),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(0.625),to_float(0.625),to_float(0.250),to_float(-0.875)),
    (to_float(0.250),to_float(-0.875),to_float(0.625),to_float(0.000),to_float(-0.875),to_float(-0.125),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(-0.500),to_float(-0.750),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(0.500),to_float(-0.125),to_float(0.125),to_float(-0.125)),
    (to_float(0.500),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(0.625),to_float(-0.625),to_float(0.875),to_float(-0.125),to_float(-0.750),to_float(0.875),to_float(-0.625),to_float(0.500),to_float(-0.125),to_float(0.500),to_float(-0.875),to_float(0.000),to_float(0.375),to_float(-0.875)),
    (to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(-0.375),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(0.750),to_float(0.875),to_float(0.250),to_float(0.625),to_float(0.125),to_float(0.750),to_float(-0.375),to_float(0.875),to_float(0.500),to_float(-0.875)),
    (to_float(-0.250),to_float(-0.875),to_float(0.375),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(0.500),to_float(0.125),to_float(0.750),to_float(0.625),to_float(-0.375),to_float(-0.875),to_float(0.625),to_float(0.750),to_float(-0.875)),
    (to_float(0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.000),to_float(0.750),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(-0.250),to_float(-0.875),to_float(-0.625),to_float(0.625),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(-0.875),to_float(-0.750),to_float(0.250),to_float(0.250),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(0.000)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.875),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.875),to_float(-0.250),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.250),to_float(-0.875)),
    (to_float(0.750),to_float(-0.875),to_float(0.125),to_float(-0.250),to_float(0.000),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(-0.750),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875)),
    (to_float(0.625),to_float(0.250),to_float(-0.625),to_float(-0.375),to_float(-0.125),to_float(-0.625),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.375),to_float(0.875),to_float(0.125),to_float(0.625),to_float(-0.750),to_float(-0.375),to_float(-0.375)),
    (to_float(-0.375),to_float(0.875),to_float(-0.625),to_float(-0.375),to_float(0.125),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.375),to_float(-0.875),to_float(0.000),to_float(-0.250),to_float(0.750),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(-0.625),to_float(0.125),to_float(-0.125)),
    (to_float(-0.500),to_float(0.125),to_float(0.750),to_float(0.875),to_float(-0.625),to_float(0.000),to_float(-0.375),to_float(-0.500),to_float(0.750),to_float(0.375),to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.000),to_float(-0.625),to_float(-0.250),to_float(0.125),to_float(-0.125)),
    (to_float(-0.250),to_float(-0.375),to_float(0.500),to_float(-0.250),to_float(0.625),to_float(0.000),to_float(-0.125),to_float(0.875),to_float(0.000),to_float(0.500),to_float(-0.125),to_float(-0.500),to_float(0.000),to_float(0.250),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(-0.500),to_float(0.250),to_float(0.000)),
    (to_float(0.375),to_float(0.375),to_float(0.625),to_float(0.500),to_float(-0.500),to_float(0.375),to_float(0.250),to_float(-0.750),to_float(0.375),to_float(0.750),to_float(0.000),to_float(0.375),to_float(-0.125),to_float(-0.250),to_float(-0.750),to_float(0.000),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(-0.250),to_float(0.125),to_float(-0.375),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(0.375),to_float(-0.250),to_float(0.625),to_float(0.500),to_float(-0.625),to_float(-0.500),to_float(0.375)),
    (to_float(0.250),to_float(-0.250),to_float(-0.250),to_float(0.000),to_float(-0.250),to_float(0.625),to_float(0.625),to_float(-0.500),to_float(0.000),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.500),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.500)),
    (to_float(-0.250),to_float(0.500),to_float(0.375),to_float(-0.375),to_float(0.500),to_float(0.875),to_float(-0.375),to_float(0.000),to_float(0.375),to_float(0.250),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.250),to_float(0.625),to_float(0.250),to_float(-0.125),to_float(-0.500),to_float(-0.125),to_float(-0.125)),
    (to_float(0.375),to_float(-0.125),to_float(0.250),to_float(0.125),to_float(0.000),to_float(0.500),to_float(0.125),to_float(0.250),to_float(0.875),to_float(-0.750),to_float(0.375),to_float(0.250),to_float(0.125),to_float(-0.500),to_float(0.625),to_float(-0.125),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(-0.125)),
    (to_float(0.500),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.500),to_float(0.250),to_float(0.125),to_float(0.125),to_float(0.625),to_float(0.250),to_float(-0.375),to_float(-0.125),to_float(0.125),to_float(0.500),to_float(-0.250),to_float(0.125),to_float(0.000),to_float(-0.750),to_float(0.000),to_float(0.125)),
    (to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.500),to_float(0.125),to_float(-0.125),to_float(-0.750),to_float(0.000),to_float(0.875),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.375),to_float(-0.500),to_float(-0.375),to_float(-0.500),to_float(-0.125),to_float(-0.250)),
    (to_float(0.250),to_float(0.250),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(0.500),to_float(0.000),to_float(-0.500),to_float(0.375),to_float(-0.625),to_float(-0.125),to_float(0.000),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(-0.625),to_float(-0.250),to_float(0.000)),
    (to_float(0.250),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.875),to_float(0.375),to_float(0.000),to_float(-0.500),to_float(0.375),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.375),to_float(0.250),to_float(0.500),to_float(0.375),to_float(-0.750),to_float(-0.125),to_float(-0.250)),
    (to_float(0.000),to_float(0.000),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(-0.750),to_float(0.250),to_float(-0.375),to_float(0.250),to_float(0.250),to_float(0.000),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(-0.625),to_float(-0.500),to_float(-0.125),to_float(-0.500)),
    (to_float(0.250),to_float(0.250),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(0.250),to_float(-0.500),to_float(0.375),to_float(-0.125),to_float(-0.375),to_float(0.250),to_float(0.000),to_float(0.125),to_float(-0.875),to_float(-0.375),to_float(-0.250),to_float(-0.875),to_float(-0.500),to_float(-0.750)),
    (to_float(-0.125),to_float(-0.375),to_float(-0.250),to_float(0.625),to_float(-0.875),to_float(0.000),to_float(-0.250),to_float(-0.375),to_float(-0.625),to_float(0.250),to_float(0.000),to_float(0.625),to_float(0.500),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(-0.500),to_float(0.000)),
    (to_float(-0.375),to_float(-0.750),to_float(-0.250),to_float(0.375),to_float(-0.875),to_float(0.500),to_float(0.375),to_float(-0.500),to_float(0.500),to_float(-0.375),to_float(-0.625),to_float(0.125),to_float(0.750),to_float(0.625),to_float(-0.750),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(0.000),to_float(-0.875)),
    (to_float(-0.125),to_float(-0.625),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(-0.625),to_float(0.750),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(-0.625),to_float(0.250),to_float(0.875),to_float(-0.625),to_float(-0.250),to_float(-0.875)),
    (to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(-0.375),to_float(0.750),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.125)),
    (to_float(0.875),to_float(0.000),to_float(-0.875),to_float(0.000),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(-0.625),to_float(0.625),to_float(-0.250),to_float(0.875),to_float(0.625),to_float(-0.125),to_float(0.250),to_float(-0.875),to_float(0.000),to_float(0.500),to_float(-0.625)),
    (to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(-0.375),to_float(-0.625),to_float(0.875),to_float(0.375),to_float(0.000),to_float(0.250),to_float(0.000),to_float(0.875),to_float(0.750),to_float(-0.875)),
    (to_float(0.625),to_float(-0.875),to_float(0.500),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(0.625),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.750),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(0.375),to_float(0.250),to_float(0.875),to_float(-0.875)),
    (to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(-0.250),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(0.750),to_float(0.375)),
    (to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125)),
    (to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.500),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(0.625),to_float(-0.625),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(-0.625),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(-0.375)),
    (to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(-0.375),to_float(0.500),to_float(-0.250),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.625),to_float(-0.125),to_float(0.250),to_float(-0.625),to_float(-0.625),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.125)),
    (to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(-0.500),to_float(0.875),to_float(0.375),to_float(0.000),to_float(-0.500),to_float(0.750),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(-0.250)),
    (to_float(-0.875),to_float(0.500),to_float(0.500),to_float(0.875),to_float(0.250),to_float(0.750),to_float(-0.125),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.375),to_float(-0.500),to_float(0.125),to_float(-0.875),to_float(0.250),to_float(-0.250),to_float(-0.125)),
    (to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.250),to_float(0.125),to_float(0.250),to_float(0.125),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(0.500),to_float(0.375),to_float(-0.875),to_float(0.375),to_float(-0.625),to_float(0.000)),
    (to_float(-0.125),to_float(0.250),to_float(0.250),to_float(-0.250),to_float(0.250),to_float(0.000),to_float(0.375),to_float(0.000),to_float(-0.125),to_float(0.875),to_float(0.000),to_float(0.125),to_float(-0.250),to_float(-0.250),to_float(-0.375),to_float(0.125),to_float(-0.500),to_float(-0.250),to_float(-0.500),to_float(0.125)),
    (to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(-0.125),to_float(-0.750),to_float(0.000),to_float(0.500),to_float(-0.750),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(-0.125),to_float(-0.250),to_float(-0.250),to_float(0.125),to_float(0.250),to_float(0.125),to_float(-0.250),to_float(-0.375),to_float(-0.375)),
    (to_float(-0.125),to_float(-0.625),to_float(-0.500),to_float(0.375),to_float(-0.625),to_float(-0.625),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(0.625),to_float(-0.625),to_float(-0.375),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(-0.500),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.250)),
    (to_float(0.375),to_float(0.000),to_float(-0.250),to_float(-0.875),to_float(-0.125),to_float(-0.375),to_float(-0.125),to_float(0.250),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(-0.250),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(0.250),to_float(-0.625),to_float(-0.375),to_float(0.250),to_float(-0.125)),
    (to_float(0.250),to_float(-0.250),to_float(0.500),to_float(0.250),to_float(0.375),to_float(0.125),to_float(0.125),to_float(-0.750),to_float(0.375),to_float(-0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.250),to_float(0.375),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.625)),
    (to_float(-0.500),to_float(0.125),to_float(0.375),to_float(0.250),to_float(0.250),to_float(-0.750),to_float(0.375),to_float(-0.375),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.250),to_float(0.500),to_float(0.125),to_float(0.750),to_float(-0.500),to_float(0.250),to_float(0.625)),
    (to_float(0.375),to_float(0.000),to_float(-0.625),to_float(-0.750),to_float(-0.750),to_float(-0.250),to_float(0.000),to_float(-0.375),to_float(0.625),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(-0.250),to_float(0.250),to_float(0.500),to_float(0.250),to_float(-0.625),to_float(-0.125),to_float(-0.625)),
    (to_float(-0.500),to_float(0.625),to_float(0.125),to_float(0.250),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(-0.750),to_float(-0.125),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(0.000),to_float(-0.625),to_float(-0.250),to_float(-0.375),to_float(-0.375),to_float(-0.750),to_float(-0.375)),
    (to_float(0.375),to_float(-0.125),to_float(-0.375),to_float(-0.250),to_float(-0.250),to_float(0.375),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(0.250),to_float(0.000),to_float(0.125),to_float(0.375),to_float(0.375),to_float(-0.500),to_float(-0.625),to_float(-0.500),to_float(-0.250),to_float(-0.875)),
    (to_float(-0.625),to_float(-0.250),to_float(-0.750),to_float(-0.125),to_float(-0.625),to_float(-0.375),to_float(-0.375),to_float(-0.125),to_float(0.875),to_float(-0.250),to_float(-0.250),to_float(-0.625),to_float(-0.625),to_float(0.250),to_float(-0.500),to_float(0.000),to_float(-0.625),to_float(-0.625),to_float(-0.375),to_float(-0.125)),
    (to_float(0.000),to_float(0.375),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(-0.750),to_float(0.250),to_float(0.125),to_float(0.750),to_float(0.375),to_float(-0.750),to_float(-0.250),to_float(-0.125),to_float(-0.625),to_float(-0.250),to_float(0.250),to_float(0.250),to_float(-0.625),to_float(-0.625),to_float(-0.375)),
    (to_float(0.625),to_float(0.625),to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(-0.750),to_float(-0.500),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(0.750),to_float(0.625),to_float(-0.250),to_float(0.125),to_float(-0.250),to_float(0.500),to_float(-0.375),to_float(-0.625)),
    (to_float(0.125),to_float(0.250),to_float(-0.375),to_float(-0.375),to_float(-0.750),to_float(-0.875),to_float(0.375),to_float(-0.625),to_float(-0.750),to_float(0.375),to_float(0.875),to_float(0.625),to_float(0.000),to_float(-0.250),to_float(-0.625),to_float(-0.625),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(-0.750)),
    (to_float(-0.375),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.000),to_float(-0.375),to_float(0.875),to_float(0.750),to_float(-0.875),to_float(0.125),to_float(0.125),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(0.000),to_float(-0.875)),
    (to_float(0.750),to_float(0.625),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(0.625),to_float(0.625),to_float(0.875),to_float(0.500),to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(0.250),to_float(-0.750)),
    (to_float(0.250),to_float(-0.125),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(0.750),to_float(0.875),to_float(0.875),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.750),to_float(0.000)),
    (to_float(0.750),to_float(0.375),to_float(-0.875),to_float(-0.750),to_float(-0.125),to_float(-0.875),to_float(0.750),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.625),to_float(0.000),to_float(0.625),to_float(0.875),to_float(0.875),to_float(0.125),to_float(0.250),to_float(0.000),to_float(-0.500),to_float(0.250)),
    (to_float(0.000),to_float(-0.875),to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.750),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.625),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.000),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.125)),
    (to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125)),
    (to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000)),
    (to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(0.500),to_float(-0.500),to_float(0.375),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(-0.625),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(0.875),to_float(0.250),to_float(0.625)),
    (to_float(-0.375),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.625)),
    (to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.125),to_float(-0.750),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.125),to_float(-0.375),to_float(0.750),to_float(0.875),to_float(-0.500),to_float(-0.250)),
    (to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.500),to_float(0.500),to_float(0.000),to_float(-0.875)),
    (to_float(-0.500),to_float(0.625),to_float(-0.250),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(0.375),to_float(0.375),to_float(-0.375),to_float(-0.250),to_float(0.250),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.000),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(-0.500)),
    (to_float(-0.875),to_float(0.500),to_float(0.000),to_float(0.500),to_float(0.250),to_float(0.625),to_float(0.875),to_float(0.750),to_float(-0.750),to_float(0.000),to_float(-0.875),to_float(-0.250),to_float(-0.250),to_float(0.625),to_float(0.000),to_float(-0.375),to_float(-0.250),to_float(0.750),to_float(0.125),to_float(-0.750)),
    (to_float(-0.125),to_float(-0.500),to_float(-0.500),to_float(-0.500),to_float(0.375),to_float(0.250),to_float(-0.125),to_float(0.250),to_float(0.625),to_float(0.000),to_float(0.125),to_float(-0.375),to_float(0.375),to_float(0.625),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(-0.500),to_float(0.625),to_float(0.250)),
    (to_float(-0.625),to_float(-0.750),to_float(-0.875),to_float(0.375),to_float(0.000),to_float(0.375),to_float(0.875),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.375),to_float(0.000),to_float(-0.375),to_float(0.250),to_float(-0.250),to_float(0.125),to_float(-0.875),to_float(-0.250),to_float(0.625),to_float(0.375)),
    (to_float(-0.375),to_float(0.625),to_float(-0.875),to_float(-0.750),to_float(-0.375),to_float(0.875),to_float(-0.750),to_float(-0.500),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(0.750),to_float(-0.375),to_float(0.500),to_float(0.000),to_float(0.625),to_float(0.125),to_float(0.250)),
    (to_float(0.000),to_float(0.625),to_float(-0.875),to_float(-0.250),to_float(-0.375),to_float(-0.250),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.625),to_float(-0.625),to_float(0.125),to_float(0.500),to_float(0.125),to_float(0.875),to_float(-0.250),to_float(0.625)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(-0.375),to_float(0.250),to_float(0.750),to_float(0.000),to_float(0.500),to_float(0.000),to_float(-0.500),to_float(-0.750),to_float(0.125),to_float(0.625),to_float(0.250),to_float(-0.375),to_float(0.000),to_float(-0.500),to_float(0.125),to_float(0.625)),
    (to_float(0.000),to_float(-0.625),to_float(-0.875),to_float(0.625),to_float(-0.375),to_float(0.125),to_float(-0.250),to_float(-0.125),to_float(0.625),to_float(0.625),to_float(-0.625),to_float(-0.625),to_float(0.625),to_float(-0.250),to_float(0.125),to_float(0.375),to_float(0.000),to_float(0.375),to_float(-0.375),to_float(0.500)),
    (to_float(-0.625),to_float(0.250),to_float(-0.875),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.500),to_float(0.000),to_float(0.000),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(-0.250),to_float(-0.125),to_float(-0.375),to_float(-0.250),to_float(0.250),to_float(-0.500),to_float(-0.125)),
    (to_float(-0.125),to_float(0.250),to_float(-0.750),to_float(-0.250),to_float(-0.500),to_float(-0.750),to_float(0.250),to_float(0.000),to_float(-0.500),to_float(0.000),to_float(-0.375),to_float(-0.500),to_float(0.125),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(0.250),to_float(0.125),to_float(0.000),to_float(-0.750)),
    (to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.375),to_float(-0.750),to_float(0.750),to_float(-0.875),to_float(0.500),to_float(0.375),to_float(0.250),to_float(0.000),to_float(0.750),to_float(0.625),to_float(0.250),to_float(0.000),to_float(0.000),to_float(0.750),to_float(0.500),to_float(0.375)),
    (to_float(0.125),to_float(-0.500),to_float(-0.750),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.000),to_float(0.375),to_float(0.875),to_float(-0.250),to_float(0.750),to_float(0.500),to_float(0.125),to_float(0.000),to_float(0.625),to_float(-0.375)),
    (to_float(0.250),to_float(0.250),to_float(-0.875),to_float(-0.500),to_float(-0.250),to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(0.875),to_float(-0.125),to_float(0.125),to_float(-0.500),to_float(-0.125),to_float(-0.500),to_float(0.250),to_float(0.250),to_float(-0.625),to_float(0.625),to_float(0.125),to_float(-0.875)),
    (to_float(0.500),to_float(0.625),to_float(-0.875),to_float(0.500),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(0.000),to_float(0.500),to_float(-0.625),to_float(-0.875),to_float(0.000),to_float(0.375),to_float(0.375)),
    (to_float(-0.125),to_float(0.750),to_float(-0.875),to_float(0.250),to_float(0.125),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.500),to_float(-0.250),to_float(-0.750),to_float(0.000),to_float(0.250),to_float(-0.875),to_float(0.375),to_float(-0.500),to_float(-0.125)),
    (to_float(0.250),to_float(0.125),to_float(-0.875),to_float(-0.750),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.875),to_float(0.375),to_float(-0.500),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.375)),
    (to_float(0.000),to_float(-0.500),to_float(-0.875),to_float(-0.375),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(0.875),to_float(0.625),to_float(0.000),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(-0.750)),
    (to_float(0.875),to_float(0.000),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(0.750),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.500),to_float(0.000),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(0.625),to_float(0.625),to_float(0.500),to_float(-0.875)),
    (to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.625),to_float(0.875),to_float(0.250),to_float(-0.125),to_float(0.875),to_float(0.000),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.625),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(0.125)),
    (to_float(0.750),to_float(-0.875),to_float(0.000),to_float(0.750),to_float(0.125),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.250),to_float(-0.500),to_float(0.875),to_float(-0.875),to_float(0.000)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125)),
    (to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125)),
    (to_float(0.000),to_float(0.125),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(0.875),to_float(-0.500),to_float(0.250),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(-0.750),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(0.875)),
    (to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(-0.625),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.000)),
    (to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(-0.625),to_float(0.500),to_float(0.750),to_float(-0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(-0.375),to_float(-0.250),to_float(-0.875),to_float(0.250),to_float(-0.750),to_float(-0.375),to_float(0.625),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.375)),
    (to_float(0.625),to_float(-0.375),to_float(-0.875),to_float(0.625),to_float(0.375),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(-0.875),to_float(0.375),to_float(0.750),to_float(0.000),to_float(0.750),to_float(-0.875),to_float(-0.750),to_float(0.500),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(-0.250)),
    (to_float(-0.875),to_float(0.250),to_float(-0.875),to_float(0.750),to_float(0.375),to_float(0.250),to_float(0.250),to_float(-0.250),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.750),to_float(0.125),to_float(-0.875),to_float(-0.375),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125)),
    (to_float(-0.875),to_float(0.375),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.500),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(0.375),to_float(-0.125),to_float(-0.250),to_float(-0.250),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(-0.875),to_float(0.500),to_float(-0.125)),
    (to_float(-0.625),to_float(-0.125),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(-0.625),to_float(-0.375),to_float(-0.875),to_float(0.250),to_float(-0.750),to_float(0.875),to_float(0.375),to_float(-0.750),to_float(-0.875),to_float(0.250),to_float(-0.125),to_float(-0.750),to_float(0.375),to_float(0.000)),
    (to_float(0.500),to_float(0.375),to_float(-0.875),to_float(-0.375),to_float(0.500),to_float(-0.500),to_float(-0.875),to_float(-0.500),to_float(-0.250),to_float(0.250),to_float(-0.250),to_float(0.250),to_float(0.500),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(0.000),to_float(0.125),to_float(0.875),to_float(-0.125)),
    (to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.250),to_float(-0.625),to_float(0.250),to_float(0.250),to_float(-0.750),to_float(-0.500),to_float(-0.875),to_float(-0.250),to_float(0.000),to_float(-0.500),to_float(0.250),to_float(0.875),to_float(0.125)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(0.750),to_float(0.250),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(0.625),to_float(0.000),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.125),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(-0.125),to_float(0.375),to_float(-0.375),to_float(-0.875),to_float(-0.125),to_float(-0.375),to_float(0.500),to_float(-0.500),to_float(-0.375),to_float(0.000),to_float(0.625),to_float(-0.625),to_float(-0.250),to_float(0.875),to_float(0.875)),
    (to_float(-0.625),to_float(0.250),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(-0.375),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.500),to_float(0.000),to_float(0.875),to_float(0.875)),
    (to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.625),to_float(-0.375),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(-0.375),to_float(0.750),to_float(0.250),to_float(-0.750),to_float(-0.875),to_float(-0.125),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(-0.750)),
    (to_float(-0.250),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.500),to_float(0.000),to_float(-0.500),to_float(-0.875),to_float(0.000),to_float(0.000),to_float(0.500),to_float(0.125),to_float(-0.625),to_float(-0.875),to_float(-0.375),to_float(-0.375),to_float(-0.750),to_float(0.875),to_float(-0.125)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.625),to_float(0.000),to_float(0.375),to_float(-0.875),to_float(-0.250),to_float(-0.375),to_float(0.000),to_float(-0.875),to_float(0.125),to_float(0.375),to_float(0.500),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(-0.375)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.625),to_float(0.625),to_float(0.125),to_float(-0.875),to_float(0.625),to_float(-0.500),to_float(-0.250),to_float(-0.250),to_float(0.375),to_float(-0.875),to_float(-0.125),to_float(0.875),to_float(-0.375)),
    (to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.375),to_float(-0.125),to_float(0.750),to_float(-0.375),to_float(0.125),to_float(0.875),to_float(0.625),to_float(0.250),to_float(0.500),to_float(-0.875),to_float(-0.500),to_float(-0.500),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(-0.875)),
    (to_float(-0.500),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.375),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(-0.625),to_float(-0.500),to_float(0.875),to_float(0.875)),
    (to_float(-0.125),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(-0.250),to_float(-0.250),to_float(-0.875),to_float(0.625),to_float(0.875),to_float(0.625),to_float(0.875),to_float(-0.875),to_float(-0.250),to_float(0.750),to_float(-0.875),to_float(-0.125),to_float(0.375),to_float(-0.500)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.750),to_float(-0.500),to_float(-0.875),to_float(0.000),to_float(-0.375),to_float(0.000),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.375),to_float(-0.875),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.125)),
    (to_float(-0.125),to_float(-0.750),to_float(-0.500),to_float(0.500),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.250),to_float(-0.250),to_float(-0.250),to_float(0.250),to_float(-0.125),to_float(-0.875),to_float(-0.500),to_float(0.375),to_float(0.250),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(-0.125)),
    (to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000)),
    (to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(-0.625),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(-0.625),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.250),to_float(0.375),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.750),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.375),to_float(0.875),to_float(-0.375),to_float(0.125),to_float(0.625),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(-0.375),to_float(-0.125),to_float(0.875),to_float(-0.500),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.000),to_float(0.500),to_float(0.875),to_float(-0.500),to_float(0.000),to_float(0.875),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.125),to_float(0.875),to_float(-0.375),to_float(0.875),to_float(0.625)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.625),to_float(-0.875),to_float(0.625),to_float(0.000),to_float(-0.625),to_float(-0.125),to_float(0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(-0.375),to_float(0.375),to_float(0.625),to_float(0.375),to_float(0.625),to_float(0.625)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.500),to_float(-0.750),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.625),to_float(0.000),to_float(-0.875),to_float(-0.375),to_float(0.125),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.000),to_float(-0.875),to_float(0.375),to_float(0.625),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.500),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.375),to_float(-0.875),to_float(-0.375),to_float(-0.250),to_float(0.625),to_float(-0.500),to_float(-0.875),to_float(-0.250),to_float(0.125),to_float(0.875),to_float(0.750),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.625),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(0.875),to_float(-0.125),to_float(0.875),to_float(-0.250)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(0.625),to_float(-0.625),to_float(0.875),to_float(-0.875),to_float(-0.500),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.750)),
    (to_float(-0.125),to_float(0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(0.375),to_float(0.625),to_float(-0.750),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.625),to_float(0.750),to_float(-0.625),to_float(0.500),to_float(0.875),to_float(-0.125)),
    (to_float(-0.250),to_float(0.625),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.500),to_float(0.625),to_float(-0.625),to_float(-0.875),to_float(0.250),to_float(0.875),to_float(0.750),to_float(-0.750),to_float(-0.875),to_float(-0.375),to_float(0.750),to_float(0.125),to_float(0.750),to_float(0.500),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(-0.125),to_float(-0.875),to_float(-0.375),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(-0.250),to_float(0.000),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(-0.875),to_float(0.500),to_float(-0.875),to_float(-0.875),to_float(-0.500),to_float(0.875),to_float(0.875),to_float(0.500),to_float(-0.750),to_float(-0.875),to_float(0.750),to_float(0.000),to_float(0.125),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.875),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.125),to_float(-0.875),to_float(0.500),to_float(0.875),to_float(-0.125),to_float(-0.625),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.875),to_float(0.000),to_float(0.500),to_float(-0.875),to_float(-0.125),to_float(0.625),to_float(0.875),to_float(0.500),to_float(0.875),to_float(-0.875),to_float(-0.375),to_float(-0.875),to_float(0.375),to_float(0.875),to_float(0.250),to_float(0.875),to_float(-0.875),to_float(0.500)),
    (to_float(-0.750),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.500),to_float(-0.625),to_float(-0.750),to_float(-0.375),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.000),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.625)),
    (to_float(0.125),to_float(0.875),to_float(-0.875),to_float(0.875),to_float(0.375),to_float(-0.250),to_float(-0.875),to_float(-0.625),to_float(0.750),to_float(0.875),to_float(0.875),to_float(-0.125),to_float(-0.875),to_float(-0.875),to_float(-0.875),to_float(0.750),to_float(0.750),to_float(0.000),to_float(0.875),to_float(0.875)),
    (to_float(-0.875),to_float(0.875),to_float(-0.750),to_float(0.500),to_float(0.125),to_float(-0.125),to_float(0.125),to_float(0.250),to_float(-0.875),to_float(-0.875),to_float(0.875),to_float(0.125),to_float(-0.875),to_float(-0.875),to_float(-0.125),to_float(0.375),to_float(0.125),to_float(-0.875),to_float(0.875),to_float(0.875)),
    (to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.125),to_float(0.125),to_float(0.000)),
    (to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(-0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000)),
    (to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(-0.125),to_float(0.125),to_float(0.000),to_float(0.000),to_float(-0.125)),
    (to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.000),to_float(0.125)));

end mulmat_mem;