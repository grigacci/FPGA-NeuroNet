library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.bfloat_pkg.ALL;

package input_data is
    type input_array is array(natural range<>, natural range<>) of bfloat16;

    --Image of index 1 , representation of the number 2

    constant input_image : input_array(27 downto 0,27 downto 0) := 
    ((to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00000823),to_bfloat16(-0.00003058),to_bfloat16(-0.00001407),to_bfloat16(-0.00000060),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00000101),to_bfloat16(-0.00000358),to_bfloat16(-0.00003624),to_bfloat16(-0.00009483),to_bfloat16(-0.00017083),to_bfloat16(-0.00025034),to_bfloat16(-0.00046921),to_bfloat16(-0.00062799),to_bfloat16(-0.00068045),to_bfloat16(-0.00069332),to_bfloat16(-0.00073957),to_bfloat16(-0.00068045),to_bfloat16(-0.00073004),to_bfloat16(-0.00060034),to_bfloat16(-0.00039101),to_bfloat16(-0.00027823),to_bfloat16(-0.00021017),to_bfloat16(-0.00008345),to_bfloat16(-0.00003940),to_bfloat16(-0.00001383),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00000417),to_bfloat16(-0.00000274),to_bfloat16(-0.00002712),to_bfloat16(-0.00002140),to_bfloat16(-0.00018394),to_bfloat16(-0.00054073),to_bfloat16(-0.00103188),to_bfloat16(-0.00197983),to_bfloat16(-0.00338554),to_bfloat16(-0.00503922),to_bfloat16(-0.00730515),to_bfloat16(-0.00988007),to_bfloat16(-0.01250458),to_bfloat16(-0.01416016),to_bfloat16(-0.01454163),to_bfloat16(-0.01325226),to_bfloat16(-0.01094818),to_bfloat16(-0.00798798),to_bfloat16(-0.00469589),to_bfloat16(-0.00247383),to_bfloat16(-0.00115681),to_bfloat16(-0.00036716),to_bfloat16(-0.00013757),to_bfloat16(-0.00003374),to_bfloat16(0.00000000),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00001264),to_bfloat16(-0.00002283),to_bfloat16(-0.00004697),to_bfloat16(-0.00027251),to_bfloat16(-0.00082827),to_bfloat16(-0.00213242),to_bfloat16(-0.00450897),to_bfloat16(-0.00865936),to_bfloat16(0.43896484),to_bfloat16(0.46704102),to_bfloat16(0.63916016),to_bfloat16(0.95800781),to_bfloat16(0.94970703),to_bfloat16(0.53417969),to_bfloat16(0.31201172),to_bfloat16(-0.04614258),to_bfloat16(-0.03729248),to_bfloat16(-0.02680969),to_bfloat16(-0.01638794),to_bfloat16(-0.00888824),to_bfloat16(-0.00414276),to_bfloat16(-0.00161362),to_bfloat16(-0.00063324),to_bfloat16(-0.00010848),to_bfloat16(-0.00001097),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(-0.00000250),to_bfloat16(-0.00002038),to_bfloat16(-0.00005603),to_bfloat16(-0.00031590),to_bfloat16(-0.00160217),to_bfloat16(-0.00407410),to_bfloat16(-0.00945282),to_bfloat16(-0.01866150),to_bfloat16(0.62744141),to_bfloat16(0.93652344),to_bfloat16(0.91210938),to_bfloat16(0.88281250),to_bfloat16(0.85058594),to_bfloat16(0.82470703),to_bfloat16(0.81152344),to_bfloat16(0.67822266),to_bfloat16(-0.03576660),to_bfloat16(-0.12237549),to_bfloat16(-0.08953857),to_bfloat16(-0.05792236),to_bfloat16(-0.03384399),to_bfloat16(-0.01776123),to_bfloat16(-0.00834656),to_bfloat16(-0.00337029),to_bfloat16(-0.00081158),to_bfloat16(-0.00011581),to_bfloat16(-0.00000793)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00004029),to_bfloat16(-0.00024748),to_bfloat16(-0.00154495),to_bfloat16(-0.00571823),to_bfloat16(-0.01401520),to_bfloat16(-0.02822876),to_bfloat16(0.60937500),to_bfloat16(0.90527344),to_bfloat16(0.86523438),to_bfloat16(0.81542969),to_bfloat16(0.60205078),to_bfloat16(0.26635742),to_bfloat16(0.35498047),to_bfloat16(0.63427734),to_bfloat16(0.64062500),to_bfloat16(0.16333008),to_bfloat16(-0.25756836),to_bfloat16(-0.19445801),to_bfloat16(-0.13415527),to_bfloat16(-0.08404541),to_bfloat16(-0.04840088),to_bfloat16(-0.02593994),to_bfloat16(-0.01168823),to_bfloat16(-0.00329590),to_bfloat16(-0.00055313),to_bfloat16(-0.00001836)),(
to_bfloat16(0.00000000),to_bfloat16(-0.00000072),to_bfloat16(-0.00010741),to_bfloat16(-0.00086498),to_bfloat16(-0.00437164),to_bfloat16(-0.01284790),to_bfloat16(-0.02905273),to_bfloat16(0.14746094),to_bfloat16(0.88232422),to_bfloat16(0.84277344),to_bfloat16(0.61279297),to_bfloat16(-0.15209961),to_bfloat16(-0.30175781),to_bfloat16(-0.41503906),to_bfloat16(-0.43945312),to_bfloat16(0.31982422),to_bfloat16(0.51269531),to_bfloat16(0.10913086),to_bfloat16(-0.37548828),to_bfloat16(-0.29370117),to_bfloat16(-0.21105957),to_bfloat16(-0.13793945),to_bfloat16(-0.08197021),to_bfloat16(-0.04470825),to_bfloat16(-0.02104187),to_bfloat16(-0.00724792),to_bfloat16(-0.00145626),to_bfloat16(-0.00011837)),(
to_bfloat16(-0.00000304),to_bfloat16(-0.00007707),to_bfloat16(-0.00042057),to_bfloat16(-0.00232697),to_bfloat16(-0.00903320),to_bfloat16(-0.02316284),to_bfloat16(-0.04858398),to_bfloat16(0.21313477),to_bfloat16(0.83886719),to_bfloat16(0.60986328),to_bfloat16(-0.19042969),to_bfloat16(-0.36767578),to_bfloat16(-0.43579102),to_bfloat16(-0.48828125),to_bfloat16(-0.04199219),to_bfloat16(0.43994141),to_bfloat16(0.46728516),to_bfloat16(-0.24096680),to_bfloat16(-0.44360352),to_bfloat16(-0.36621094),to_bfloat16(-0.27246094),to_bfloat16(-0.18298340),to_bfloat16(-0.10992432),to_bfloat16(-0.05938721),to_bfloat16(-0.02748108),to_bfloat16(-0.01009369),to_bfloat16(-0.00200462),to_bfloat16(-0.00012457)),(
to_bfloat16(-0.00001591),to_bfloat16(-0.00019848),to_bfloat16(-0.00128651),to_bfloat16(-0.00514603),to_bfloat16(-0.01464081),to_bfloat16(-0.03314209),to_bfloat16(-0.06567383),to_bfloat16(-0.11560059),to_bfloat16(-0.06225586),to_bfloat16(-0.19580078),to_bfloat16(-0.35278320),to_bfloat16(-0.42382812),to_bfloat16(-0.46655273),to_bfloat16(-0.48193359),to_bfloat16(0.33569336),to_bfloat16(0.51074219),to_bfloat16(0.50878906),to_bfloat16(-0.22314453),to_bfloat16(-0.45410156),to_bfloat16(-0.39306641),to_bfloat16(-0.30200195),to_bfloat16(-0.20666504),to_bfloat16(-0.12426758),to_bfloat16(-0.06390381),to_bfloat16(-0.02807617),to_bfloat16(-0.01018524),to_bfloat16(-0.00188160),to_bfloat16(-0.00010616)),(
to_bfloat16(-0.00001901),to_bfloat16(-0.00031042),to_bfloat16(-0.00200081),to_bfloat16(-0.00671768),to_bfloat16(-0.01736450),to_bfloat16(-0.03829956),to_bfloat16(-0.07629395),to_bfloat16(-0.13476562),to_bfloat16(-0.21362305),to_bfloat16(-0.30517578),to_bfloat16(-0.38696289),to_bfloat16(-0.43212891),to_bfloat16(-0.43286133),to_bfloat16(0.04858398),to_bfloat16(0.57812500),to_bfloat16(0.60009766),to_bfloat16(0.36596680),to_bfloat16(-0.39404297),to_bfloat16(-0.43383789),to_bfloat16(-0.38720703),to_bfloat16(-0.30102539),to_bfloat16(-0.20593262),to_bfloat16(-0.12286377),to_bfloat16(-0.06011963),to_bfloat16(-0.02328491),to_bfloat16(-0.00741577),to_bfloat16(-0.00137424),to_bfloat16(-0.00011021)),(
to_bfloat16(-0.00002605),to_bfloat16(-0.00038505),to_bfloat16(-0.00204277),to_bfloat16(-0.00654221),to_bfloat16(-0.01675415),to_bfloat16(-0.03857422),to_bfloat16(-0.08026123),to_bfloat16(-0.14526367),to_bfloat16(-0.23327637),to_bfloat16(-0.32568359),to_bfloat16(-0.39160156),to_bfloat16(-0.40307617),to_bfloat16(-0.06982422),to_bfloat16(0.64062500),to_bfloat16(0.67773438),to_bfloat16(0.57226562),to_bfloat16(-0.12060547),to_bfloat16(-0.40795898),to_bfloat16(-0.41503906),to_bfloat16(-0.36816406),to_bfloat16(-0.28076172),to_bfloat16(-0.18872070),to_bfloat16(-0.11126709),to_bfloat16(-0.05273438),to_bfloat16(-0.01797485),to_bfloat16(-0.00449371),to_bfloat16(-0.00086641),to_bfloat16(-0.00007319)),(
to_bfloat16(-0.00002319),to_bfloat16(-0.00029850),to_bfloat16(-0.00164413),to_bfloat16(-0.00500107),to_bfloat16(-0.01424408),to_bfloat16(-0.03732300),to_bfloat16(-0.08258057),to_bfloat16(-0.15563965),to_bfloat16(-0.25024414),to_bfloat16(-0.34057617),to_bfloat16(-0.38574219),to_bfloat16(-0.37060547),to_bfloat16(0.18090820),to_bfloat16(0.70214844),to_bfloat16(0.69091797),to_bfloat16(0.22875977),to_bfloat16(-0.38012695),to_bfloat16(-0.41992188),to_bfloat16(-0.41210938),to_bfloat16(-0.34765625),to_bfloat16(-0.25366211),to_bfloat16(-0.16601562),to_bfloat16(-0.09899902),to_bfloat16(-0.04913330),to_bfloat16(-0.01558685),to_bfloat16(-0.00236130),to_bfloat16(-0.00048637),to_bfloat16(-0.00003189)),(
to_bfloat16(-0.00001484),to_bfloat16(-0.00017059),to_bfloat16(-0.00094557),to_bfloat16(-0.00343323),to_bfloat16(-0.01198578),to_bfloat16(-0.03753662),to_bfloat16(-0.08898926),to_bfloat16(-0.17016602),to_bfloat16(-0.26953125),to_bfloat16(-0.35253906),to_bfloat16(-0.38232422),to_bfloat16(0.33178711),to_bfloat16(0.64941406),to_bfloat16(0.67822266),to_bfloat16(0.27221680),to_bfloat16(-0.35034180),to_bfloat16(-0.44165039),to_bfloat16(-0.45922852),to_bfloat16(-0.41967773),to_bfloat16(-0.33007812),to_bfloat16(-0.22888184),to_bfloat16(-0.14941406),to_bfloat16(-0.09271240),to_bfloat16(-0.04965210),to_bfloat16(-0.01676941),to_bfloat16(-0.00173187),to_bfloat16(-0.00031161),to_bfloat16(-0.00003970)),(
to_bfloat16(-0.00000209),to_bfloat16(-0.00007129),to_bfloat16(-0.00047898),to_bfloat16(-0.00237274),to_bfloat16(-0.01139832),to_bfloat16(-0.04153442),to_bfloat16(-0.09979248),to_bfloat16(-0.18591309),to_bfloat16(-0.28369141),to_bfloat16(-0.35815430),to_bfloat16(-0.28076172),to_bfloat16(0.55810547),to_bfloat16(0.64892578),to_bfloat16(0.53125000),to_bfloat16(-0.29833984),to_bfloat16(-0.48437500),to_bfloat16(-0.50683594),to_bfloat16(-0.49462891),to_bfloat16(-0.42529297),to_bfloat16(-0.31713867),to_bfloat16(-0.21569824),to_bfloat16(-0.14538574),to_bfloat16(-0.09362793),to_bfloat16(-0.05328369),to_bfloat16(-0.01992798),to_bfloat16(-0.00228310),to_bfloat16(-0.00032425),to_bfloat16(-0.00004244)),(
to_bfloat16(-0.00000733),to_bfloat16(-0.00003225),to_bfloat16(-0.00021160),to_bfloat16(-0.00182056),to_bfloat16(-0.01197815),to_bfloat16(-0.04824829),to_bfloat16(-0.11145020),to_bfloat16(-0.19726562),to_bfloat16(-0.28808594),to_bfloat16(-0.35302734),to_bfloat16(0.40209961),to_bfloat16(0.62402344),to_bfloat16(0.60644531),to_bfloat16(0.09985352),to_bfloat16(-0.50878906),to_bfloat16(-0.54492188),to_bfloat16(-0.53564453),to_bfloat16(-0.50048828),to_bfloat16(-0.41796875),to_bfloat16(-0.31079102),to_bfloat16(-0.21911621),to_bfloat16(-0.15209961),to_bfloat16(-0.09973145),to_bfloat16(-0.05709839),to_bfloat16(-0.02235413),to_bfloat16(-0.00320435),to_bfloat16(-0.00036120),to_bfloat16(-0.00000864)),(
to_bfloat16(-0.00000286),to_bfloat16(-0.00001508),to_bfloat16(-0.00017619),to_bfloat16(-0.00197411),to_bfloat16(-0.01390839),to_bfloat16(-0.05627441),to_bfloat16(-0.12103271),to_bfloat16(-0.20007324),to_bfloat16(-0.27905273),to_bfloat16(-0.03027344),to_bfloat16(0.61181641),to_bfloat16(0.62011719),to_bfloat16(0.32788086),to_bfloat16(-0.43432617),to_bfloat16(-0.53027344),to_bfloat16(-0.54345703),to_bfloat16(-0.51464844),to_bfloat16(-0.47436523),to_bfloat16(-0.39575195),to_bfloat16(-0.30615234),to_bfloat16(-0.22766113),to_bfloat16(-0.16113281),to_bfloat16(-0.10540771),to_bfloat16(-0.05816650),to_bfloat16(-0.02276611),to_bfloat16(-0.00421524),to_bfloat16(-0.00057888),to_bfloat16(-0.00004232)),(
to_bfloat16(-0.00000262),to_bfloat16(-0.00001550),to_bfloat16(-0.00029039),to_bfloat16(-0.00243378),to_bfloat16(-0.01745605),to_bfloat16(-0.06457520),to_bfloat16(-0.12719727),to_bfloat16(-0.19506836),to_bfloat16(-0.18481445),to_bfloat16(0.47705078),to_bfloat16(0.66113281),to_bfloat16(0.63867188),to_bfloat16(0.15576172),to_bfloat16(-0.45263672),to_bfloat16(-0.49414062),to_bfloat16(-0.49780273),to_bfloat16(-0.47290039),to_bfloat16(-0.43432617),to_bfloat16(-0.37255859),to_bfloat16(-0.30224609),to_bfloat16(-0.23278809),to_bfloat16(-0.16418457),to_bfloat16(-0.10443115),to_bfloat16(-0.05563354),to_bfloat16(-0.02194214),to_bfloat16(-0.00502777),to_bfloat16(-0.00074816),to_bfloat16(-0.00004804)),(
to_bfloat16(0.00000000),to_bfloat16(-0.00002843),to_bfloat16(-0.00043821),to_bfloat16(-0.00372314),to_bfloat16(-0.02325439),to_bfloat16(-0.07238770),to_bfloat16(-0.13061523),to_bfloat16(-0.18823242),to_bfloat16(0.28710938),to_bfloat16(0.71777344),to_bfloat16(0.69628906),to_bfloat16(0.36035156),to_bfloat16(-0.30297852),to_bfloat16(-0.39819336),to_bfloat16(-0.43994141),to_bfloat16(-0.45092773),to_bfloat16(-0.43847656),to_bfloat16(-0.40820312),to_bfloat16(-0.36181641),to_bfloat16(-0.30175781),to_bfloat16(-0.23181152),to_bfloat16(-0.15942383),to_bfloat16(-0.09741211),to_bfloat16(-0.05014038),to_bfloat16(-0.02014160),to_bfloat16(-0.00553513),to_bfloat16(-0.00082064),to_bfloat16(-0.00003469)),(
to_bfloat16(-0.00000745),to_bfloat16(-0.00002074),to_bfloat16(-0.00070524),to_bfloat16(-0.00593948),to_bfloat16(-0.02976990),to_bfloat16(-0.07977295),to_bfloat16(-0.13635254),to_bfloat16(-0.18823242),to_bfloat16(0.74121094),to_bfloat16(0.73046875),to_bfloat16(0.70800781),to_bfloat16(-0.20141602),to_bfloat16(-0.32470703),to_bfloat16(-0.37158203),to_bfloat16(-0.41625977),to_bfloat16(-0.43823242),to_bfloat16(-0.43505859),to_bfloat16(-0.41015625),to_bfloat16(-0.36572266),to_bfloat16(-0.29931641),to_bfloat16(-0.22143555),to_bfloat16(-0.14746094),to_bfloat16(-0.08807373),to_bfloat16(-0.04446411),to_bfloat16(-0.01788330),to_bfloat16(-0.00507355),to_bfloat16(-0.00060129),to_bfloat16(-0.00004756)),(
to_bfloat16(-0.00000095),to_bfloat16(-0.00004756),to_bfloat16(-0.00111866),to_bfloat16(-0.00798035),to_bfloat16(-0.03408813),to_bfloat16(-0.08489990),to_bfloat16(-0.14392090),to_bfloat16(-0.19909668),to_bfloat16(0.72509766),to_bfloat16(0.70996094),to_bfloat16(0.68408203),to_bfloat16(-0.15478516),to_bfloat16(-0.27319336),to_bfloat16(-0.31811523),to_bfloat16(-0.36108398),to_bfloat16(-0.38208008),to_bfloat16(-0.43334961),to_bfloat16(-0.41967773),to_bfloat16(-0.34082031),to_bfloat16(-0.20263672),to_bfloat16(-0.12036133),to_bfloat16(0.01684570),to_bfloat16(0.51269531),to_bfloat16(0.55029297),to_bfloat16(0.57177734),to_bfloat16(0.56982422),to_bfloat16(0.03848267),to_bfloat16(-0.00002670)),(
to_bfloat16(0.00000000),to_bfloat16(-0.00005966),to_bfloat16(-0.00129700),to_bfloat16(-0.00881195),to_bfloat16(-0.03326416),to_bfloat16(-0.08081055),to_bfloat16(-0.14489746),to_bfloat16(-0.21008301),to_bfloat16(0.69970703),to_bfloat16(0.67089844),to_bfloat16(0.63525391),to_bfloat16(0.60595703),to_bfloat16(0.57128906),to_bfloat16(0.53027344),to_bfloat16(0.50000000),to_bfloat16(0.49780273),to_bfloat16(0.19458008),to_bfloat16(0.15307617),to_bfloat16(0.32080078),to_bfloat16(0.74902344),to_bfloat16(0.82812500),to_bfloat16(0.89062500),to_bfloat16(0.93505859),to_bfloat16(0.96289062),to_bfloat16(0.97753906),to_bfloat16(0.98535156),to_bfloat16(0.47998047),to_bfloat16(-0.00000656)),(
to_bfloat16(-0.00000209),to_bfloat16(-0.00004959),to_bfloat16(-0.00111008),to_bfloat16(-0.00718307),to_bfloat16(-0.02590942),to_bfloat16(-0.06604004),to_bfloat16(-0.12817383),to_bfloat16(-0.20141602),to_bfloat16(0.40454102),to_bfloat16(0.64746094),to_bfloat16(0.59375000),to_bfloat16(0.54882812),to_bfloat16(0.50927734),to_bfloat16(0.47900391),to_bfloat16(0.47314453),to_bfloat16(0.50048828),to_bfloat16(0.55859375),to_bfloat16(0.63867188),to_bfloat16(0.72851562),to_bfloat16(0.81005859),to_bfloat16(0.86132812),to_bfloat16(0.90136719),to_bfloat16(0.93164062),to_bfloat16(0.64404297),to_bfloat16(0.45043945),to_bfloat16(0.45532227),to_bfloat16(0.22241211),to_bfloat16(-0.00000256)),(
to_bfloat16(-0.00000203),to_bfloat16(-0.00000381),to_bfloat16(-0.00073099),to_bfloat16(-0.00424957),to_bfloat16(-0.01541138),to_bfloat16(-0.04235840),to_bfloat16(-0.09136963),to_bfloat16(-0.15869141),to_bfloat16(-0.23815918),to_bfloat16(0.14453125),to_bfloat16(0.09326172),to_bfloat16(0.03857422),to_bfloat16(0.00195312),to_bfloat16(0.15893555),to_bfloat16(0.51708984),to_bfloat16(0.56933594),to_bfloat16(0.64550781),to_bfloat16(0.34765625),to_bfloat16(0.30322266),to_bfloat16(0.36816406),to_bfloat16(0.09411621),to_bfloat16(-0.03579712),to_bfloat16(-0.01838684),to_bfloat16(-0.00868988),to_bfloat16(-0.00326157),to_bfloat16(-0.00073862),to_bfloat16(-0.00006968),to_bfloat16(-0.00000471)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00025058),to_bfloat16(-0.00163555),to_bfloat16(-0.00676727),to_bfloat16(-0.01959229),to_bfloat16(-0.04699707),to_bfloat16(-0.09350586),to_bfloat16(-0.15722656),to_bfloat16(-0.23010254),to_bfloat16(-0.30175781),to_bfloat16(-0.35961914),to_bfloat16(-0.38940430),to_bfloat16(-0.38745117),to_bfloat16(-0.35375977),to_bfloat16(-0.29516602),to_bfloat16(-0.22497559),to_bfloat16(-0.15698242),to_bfloat16(-0.09960938),to_bfloat16(-0.05953979),to_bfloat16(-0.03329468),to_bfloat16(-0.01725769),to_bfloat16(-0.00861359),to_bfloat16(-0.00383377),to_bfloat16(-0.00121212),to_bfloat16(-0.00022638),to_bfloat16(-0.00003755),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00006193),to_bfloat16(-0.00047731),to_bfloat16(-0.00212288),to_bfloat16(-0.00625229),to_bfloat16(-0.01641846),to_bfloat16(-0.03570557),to_bfloat16(-0.06573486),to_bfloat16(-0.10577393),to_bfloat16(-0.14880371),to_bfloat16(-0.18371582),to_bfloat16(-0.20153809),to_bfloat16(-0.19909668),to_bfloat16(-0.17749023),to_bfloat16(-0.14355469),to_bfloat16(-0.10717773),to_bfloat16(-0.07464600),to_bfloat16(-0.04733276),to_bfloat16(-0.02818298),to_bfloat16(-0.01546478),to_bfloat16(-0.00778580),to_bfloat16(-0.00371552),to_bfloat16(-0.00156116),to_bfloat16(-0.00039768),to_bfloat16(-0.00008667),to_bfloat16(-0.00000757),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00000614),to_bfloat16(-0.00006944),to_bfloat16(-0.00049925),to_bfloat16(-0.00185394),to_bfloat16(-0.00548935),to_bfloat16(-0.01242828),to_bfloat16(-0.02400208),to_bfloat16(-0.03839111),to_bfloat16(-0.05416870),to_bfloat16(-0.06530762),to_bfloat16(-0.07067871),to_bfloat16(-0.06945801),to_bfloat16(-0.06173706),to_bfloat16(-0.05126953),to_bfloat16(-0.04101562),to_bfloat16(-0.03044128),to_bfloat16(-0.02040100),to_bfloat16(-0.01235199),to_bfloat16(-0.00660706),to_bfloat16(-0.00322342),to_bfloat16(-0.00144768),to_bfloat16(-0.00054598),to_bfloat16(-0.00012219),to_bfloat16(-0.00001395),to_bfloat16(-0.00000679),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00000250),to_bfloat16(-0.00013852),to_bfloat16(-0.00063705),to_bfloat16(-0.00210190),to_bfloat16(-0.00468445),to_bfloat16(-0.00904846),to_bfloat16(-0.01371765),to_bfloat16(-0.01895142),to_bfloat16(-0.02336121),to_bfloat16(-0.02517700),to_bfloat16(-0.02444458),to_bfloat16(-0.02175903),to_bfloat16(-0.01737976),to_bfloat16(-0.01380920),to_bfloat16(-0.01012421),to_bfloat16(-0.00664520),to_bfloat16(-0.00394058),to_bfloat16(-0.00211143),to_bfloat16(-0.00093126),to_bfloat16(-0.00029397),to_bfloat16(-0.00006312),to_bfloat16(-0.00000203),to_bfloat16(-0.00000381),to_bfloat16(0.00000000),to_bfloat16(0.00000000)),(
to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(-0.00000989),to_bfloat16(-0.00006086),to_bfloat16(-0.00016260),to_bfloat16(-0.00034833),to_bfloat16(-0.00050068),to_bfloat16(-0.00076866),to_bfloat16(-0.00131226),to_bfloat16(-0.00167942),to_bfloat16(-0.00205421),to_bfloat16(-0.00230789),to_bfloat16(-0.00268745),to_bfloat16(-0.00231361),to_bfloat16(-0.00188541),to_bfloat16(-0.00134182),to_bfloat16(-0.00078297),to_bfloat16(-0.00034714),to_bfloat16(-0.00017822),to_bfloat16(-0.00007534),to_bfloat16(-0.00005907),to_bfloat16(-0.00000781),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000),to_bfloat16(0.00000000)));

end package;    